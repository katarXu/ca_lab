
module mem #(                   // 
    parameter  ADDR_LEN  = 11   // 
) (
    input  clk, rst,
    input  [ADDR_LEN-1:0] addr, // memory address
    output reg [31:0] rd_data,  // data read out
    input  wr_req,
    input  [31:0] wr_data       // data write in
);
localparam MEM_SIZE = 2000;
reg [31:0] ram_cell [MEM_SIZE];

always @ (posedge clk or posedge rst)
    if(rst)
        rd_data <= 0;
    else
        rd_data <= ram_cell[addr];

always @ (posedge clk)
    if(wr_req) 
        ram_cell[addr] <= wr_data;

initial begin
    // dst matrix C
    ram_cell[       0] = 32'h0;  // 32'h7906ccdf;
    ram_cell[       1] = 32'h0;  // 32'h96a700dd;
    ram_cell[       2] = 32'h0;  // 32'h3cf46b0e;
    ram_cell[       3] = 32'h0;  // 32'h261b0194;
    ram_cell[       4] = 32'h0;  // 32'he2d7c798;
    ram_cell[       5] = 32'h0;  // 32'h854d152b;
    ram_cell[       6] = 32'h0;  // 32'h19defb1a;
    ram_cell[       7] = 32'h0;  // 32'h2af51316;
    ram_cell[       8] = 32'h0;  // 32'h02f5f0f1;
    ram_cell[       9] = 32'h0;  // 32'hd8490bbb;
    ram_cell[      10] = 32'h0;  // 32'ha98bbe5d;
    ram_cell[      11] = 32'h0;  // 32'hdf955b01;
    ram_cell[      12] = 32'h0;  // 32'h56fb14bc;
    ram_cell[      13] = 32'h0;  // 32'h77daf27e;
    ram_cell[      14] = 32'h0;  // 32'h3b36e675;
    ram_cell[      15] = 32'h0;  // 32'h47eac43c;
    ram_cell[      16] = 32'h0;  // 32'hcc5b05e6;
    ram_cell[      17] = 32'h0;  // 32'hc64814eb;
    ram_cell[      18] = 32'h0;  // 32'h20be3fc9;
    ram_cell[      19] = 32'h0;  // 32'h89b83c73;
    ram_cell[      20] = 32'h0;  // 32'h00fa1ab0;
    ram_cell[      21] = 32'h0;  // 32'h21ca1d93;
    ram_cell[      22] = 32'h0;  // 32'h16758987;
    ram_cell[      23] = 32'h0;  // 32'hde7e7031;
    ram_cell[      24] = 32'h0;  // 32'hb15aa0d4;
    ram_cell[      25] = 32'h0;  // 32'h9c9a183f;
    ram_cell[      26] = 32'h0;  // 32'hcc7fa28f;
    ram_cell[      27] = 32'h0;  // 32'h5b76cdfe;
    ram_cell[      28] = 32'h0;  // 32'hfe0edfb3;
    ram_cell[      29] = 32'h0;  // 32'h4070276b;
    ram_cell[      30] = 32'h0;  // 32'hb3814d0a;
    ram_cell[      31] = 32'h0;  // 32'hcbe5a6e2;
    ram_cell[      32] = 32'h0;  // 32'h9d0115ee;
    ram_cell[      33] = 32'h0;  // 32'h7e51a635;
    ram_cell[      34] = 32'h0;  // 32'h4af98c12;
    ram_cell[      35] = 32'h0;  // 32'h94ecfb5e;
    ram_cell[      36] = 32'h0;  // 32'hd4e32e2f;
    ram_cell[      37] = 32'h0;  // 32'h574fc0de;
    ram_cell[      38] = 32'h0;  // 32'h07413ef2;
    ram_cell[      39] = 32'h0;  // 32'h6e750336;
    ram_cell[      40] = 32'h0;  // 32'hcd17e1db;
    ram_cell[      41] = 32'h0;  // 32'h73e342af;
    ram_cell[      42] = 32'h0;  // 32'h0d3cf7bc;
    ram_cell[      43] = 32'h0;  // 32'hb49d1097;
    ram_cell[      44] = 32'h0;  // 32'h56e44b32;
    ram_cell[      45] = 32'h0;  // 32'hcd3cc679;
    ram_cell[      46] = 32'h0;  // 32'h1417575e;
    ram_cell[      47] = 32'h0;  // 32'h10cfd055;
    ram_cell[      48] = 32'h0;  // 32'h587d1297;
    ram_cell[      49] = 32'h0;  // 32'h9d223789;
    ram_cell[      50] = 32'h0;  // 32'hae3aaf4e;
    ram_cell[      51] = 32'h0;  // 32'hb2b9b51d;
    ram_cell[      52] = 32'h0;  // 32'h17cdffbd;
    ram_cell[      53] = 32'h0;  // 32'hfdd9c263;
    ram_cell[      54] = 32'h0;  // 32'hd712b004;
    ram_cell[      55] = 32'h0;  // 32'h8ab30f00;
    ram_cell[      56] = 32'h0;  // 32'h5ba0b255;
    ram_cell[      57] = 32'h0;  // 32'h50298d33;
    ram_cell[      58] = 32'h0;  // 32'hcb428f5c;
    ram_cell[      59] = 32'h0;  // 32'hb66f73f8;
    ram_cell[      60] = 32'h0;  // 32'h0b2016c0;
    ram_cell[      61] = 32'h0;  // 32'h09fdc227;
    ram_cell[      62] = 32'h0;  // 32'h72efe5c4;
    ram_cell[      63] = 32'h0;  // 32'h1f46d081;
    ram_cell[      64] = 32'h0;  // 32'h839c8838;
    ram_cell[      65] = 32'h0;  // 32'hf95e6e4b;
    ram_cell[      66] = 32'h0;  // 32'hcf61d2cc;
    ram_cell[      67] = 32'h0;  // 32'he87e1ad8;
    ram_cell[      68] = 32'h0;  // 32'hcf26388c;
    ram_cell[      69] = 32'h0;  // 32'h6f7097e4;
    ram_cell[      70] = 32'h0;  // 32'h0aa9fdd0;
    ram_cell[      71] = 32'h0;  // 32'hed2dfc01;
    ram_cell[      72] = 32'h0;  // 32'h09026542;
    ram_cell[      73] = 32'h0;  // 32'h2ecb23f7;
    ram_cell[      74] = 32'h0;  // 32'hf79339a2;
    ram_cell[      75] = 32'h0;  // 32'h4f9859e9;
    ram_cell[      76] = 32'h0;  // 32'h789efc08;
    ram_cell[      77] = 32'h0;  // 32'h8de622b2;
    ram_cell[      78] = 32'h0;  // 32'h73fbe88c;
    ram_cell[      79] = 32'h0;  // 32'h97825550;
    ram_cell[      80] = 32'h0;  // 32'h61eeeb2f;
    ram_cell[      81] = 32'h0;  // 32'h0d34d015;
    ram_cell[      82] = 32'h0;  // 32'hdccf1b47;
    ram_cell[      83] = 32'h0;  // 32'ha2742fb6;
    ram_cell[      84] = 32'h0;  // 32'h787fcf67;
    ram_cell[      85] = 32'h0;  // 32'h413df402;
    ram_cell[      86] = 32'h0;  // 32'ha5a4d436;
    ram_cell[      87] = 32'h0;  // 32'hc684862d;
    ram_cell[      88] = 32'h0;  // 32'haa81c564;
    ram_cell[      89] = 32'h0;  // 32'ha4ebf34c;
    ram_cell[      90] = 32'h0;  // 32'h51ab22d4;
    ram_cell[      91] = 32'h0;  // 32'h93845c11;
    ram_cell[      92] = 32'h0;  // 32'h69b88a5f;
    ram_cell[      93] = 32'h0;  // 32'h327d623f;
    ram_cell[      94] = 32'h0;  // 32'h0939e1fe;
    ram_cell[      95] = 32'h0;  // 32'h9b03c5af;
    ram_cell[      96] = 32'h0;  // 32'hd96c6ebc;
    ram_cell[      97] = 32'h0;  // 32'h6d59bd6c;
    ram_cell[      98] = 32'h0;  // 32'hd5823a42;
    ram_cell[      99] = 32'h0;  // 32'h79ddb056;
    ram_cell[     100] = 32'h0;  // 32'hb0e90201;
    ram_cell[     101] = 32'h0;  // 32'h4c2ddfe1;
    ram_cell[     102] = 32'h0;  // 32'h92c0a757;
    ram_cell[     103] = 32'h0;  // 32'h78d9ede5;
    ram_cell[     104] = 32'h0;  // 32'hc3c90554;
    ram_cell[     105] = 32'h0;  // 32'h2978b5c4;
    ram_cell[     106] = 32'h0;  // 32'h2b3053e7;
    ram_cell[     107] = 32'h0;  // 32'h3589e59e;
    ram_cell[     108] = 32'h0;  // 32'hb4538f04;
    ram_cell[     109] = 32'h0;  // 32'h37fff18d;
    ram_cell[     110] = 32'h0;  // 32'hce4a3463;
    ram_cell[     111] = 32'h0;  // 32'h5d6600a5;
    ram_cell[     112] = 32'h0;  // 32'h17abdbae;
    ram_cell[     113] = 32'h0;  // 32'hcb799fbd;
    ram_cell[     114] = 32'h0;  // 32'h66d5b6bc;
    ram_cell[     115] = 32'h0;  // 32'h5f3805eb;
    ram_cell[     116] = 32'h0;  // 32'hf1f22a6a;
    ram_cell[     117] = 32'h0;  // 32'h5cdf02c1;
    ram_cell[     118] = 32'h0;  // 32'hd6895a25;
    ram_cell[     119] = 32'h0;  // 32'hedfb7583;
    ram_cell[     120] = 32'h0;  // 32'h74cf1bd6;
    ram_cell[     121] = 32'h0;  // 32'h9f3b7e70;
    ram_cell[     122] = 32'h0;  // 32'h1c2ca208;
    ram_cell[     123] = 32'h0;  // 32'h83a108be;
    ram_cell[     124] = 32'h0;  // 32'h1ff2e76a;
    ram_cell[     125] = 32'h0;  // 32'h21c0a546;
    ram_cell[     126] = 32'h0;  // 32'h95a290fe;
    ram_cell[     127] = 32'h0;  // 32'h256fdba3;
    ram_cell[     128] = 32'h0;  // 32'h888c74ad;
    ram_cell[     129] = 32'h0;  // 32'hc9c7b3b8;
    ram_cell[     130] = 32'h0;  // 32'hf6c1e5ff;
    ram_cell[     131] = 32'h0;  // 32'hc8f2140b;
    ram_cell[     132] = 32'h0;  // 32'hc5c8e8d9;
    ram_cell[     133] = 32'h0;  // 32'h85079be3;
    ram_cell[     134] = 32'h0;  // 32'h4961c5e8;
    ram_cell[     135] = 32'h0;  // 32'h7aaccf09;
    ram_cell[     136] = 32'h0;  // 32'h9d726659;
    ram_cell[     137] = 32'h0;  // 32'hd785fd49;
    ram_cell[     138] = 32'h0;  // 32'hbf730466;
    ram_cell[     139] = 32'h0;  // 32'h495bedee;
    ram_cell[     140] = 32'h0;  // 32'h99cfa942;
    ram_cell[     141] = 32'h0;  // 32'hc3b89225;
    ram_cell[     142] = 32'h0;  // 32'hcc075aac;
    ram_cell[     143] = 32'h0;  // 32'hb20d8ee3;
    ram_cell[     144] = 32'h0;  // 32'h72b666fa;
    ram_cell[     145] = 32'h0;  // 32'h78bf7c50;
    ram_cell[     146] = 32'h0;  // 32'h36d174e7;
    ram_cell[     147] = 32'h0;  // 32'he59119cf;
    ram_cell[     148] = 32'h0;  // 32'h423bc7ad;
    ram_cell[     149] = 32'h0;  // 32'h12c52f15;
    ram_cell[     150] = 32'h0;  // 32'h026b31df;
    ram_cell[     151] = 32'h0;  // 32'h4b1e13d2;
    ram_cell[     152] = 32'h0;  // 32'hd65f6842;
    ram_cell[     153] = 32'h0;  // 32'hdb8607a3;
    ram_cell[     154] = 32'h0;  // 32'hee196251;
    ram_cell[     155] = 32'h0;  // 32'h429c96a2;
    ram_cell[     156] = 32'h0;  // 32'hf3ca38d9;
    ram_cell[     157] = 32'h0;  // 32'h03f9d8e1;
    ram_cell[     158] = 32'h0;  // 32'h253aeb1e;
    ram_cell[     159] = 32'h0;  // 32'hb03a85e9;
    ram_cell[     160] = 32'h0;  // 32'h406a73d5;
    ram_cell[     161] = 32'h0;  // 32'h8b2b3a5b;
    ram_cell[     162] = 32'h0;  // 32'h945cd0ca;
    ram_cell[     163] = 32'h0;  // 32'hf764fdd8;
    ram_cell[     164] = 32'h0;  // 32'h5e91a26b;
    ram_cell[     165] = 32'h0;  // 32'hcc757320;
    ram_cell[     166] = 32'h0;  // 32'h73f4e06d;
    ram_cell[     167] = 32'h0;  // 32'hf578bbc7;
    ram_cell[     168] = 32'h0;  // 32'h63e8c5d8;
    ram_cell[     169] = 32'h0;  // 32'h09fa833a;
    ram_cell[     170] = 32'h0;  // 32'h7b039aeb;
    ram_cell[     171] = 32'h0;  // 32'h882ec5ce;
    ram_cell[     172] = 32'h0;  // 32'hc61f3f5e;
    ram_cell[     173] = 32'h0;  // 32'h95b501ae;
    ram_cell[     174] = 32'h0;  // 32'h91a47ee8;
    ram_cell[     175] = 32'h0;  // 32'h91251ed7;
    ram_cell[     176] = 32'h0;  // 32'h5e0e9e4c;
    ram_cell[     177] = 32'h0;  // 32'hf24af501;
    ram_cell[     178] = 32'h0;  // 32'hed95f370;
    ram_cell[     179] = 32'h0;  // 32'hb7325151;
    ram_cell[     180] = 32'h0;  // 32'h69718822;
    ram_cell[     181] = 32'h0;  // 32'h010ce755;
    ram_cell[     182] = 32'h0;  // 32'hd5c8af3e;
    ram_cell[     183] = 32'h0;  // 32'h329a1c4d;
    ram_cell[     184] = 32'h0;  // 32'hef0d85b9;
    ram_cell[     185] = 32'h0;  // 32'h84e37780;
    ram_cell[     186] = 32'h0;  // 32'h3a6563e4;
    ram_cell[     187] = 32'h0;  // 32'h47acdf88;
    ram_cell[     188] = 32'h0;  // 32'hf6fa0be8;
    ram_cell[     189] = 32'h0;  // 32'h2421fccc;
    ram_cell[     190] = 32'h0;  // 32'h883f3f07;
    ram_cell[     191] = 32'h0;  // 32'hc013edae;
    ram_cell[     192] = 32'h0;  // 32'h3190c74f;
    ram_cell[     193] = 32'h0;  // 32'hca2b75ec;
    ram_cell[     194] = 32'h0;  // 32'hb2435548;
    ram_cell[     195] = 32'h0;  // 32'h8305e7b7;
    ram_cell[     196] = 32'h0;  // 32'hd9c8bf17;
    ram_cell[     197] = 32'h0;  // 32'hfc2891b4;
    ram_cell[     198] = 32'h0;  // 32'hdedae90a;
    ram_cell[     199] = 32'h0;  // 32'h8338f57c;
    ram_cell[     200] = 32'h0;  // 32'h1c188667;
    ram_cell[     201] = 32'h0;  // 32'hde65386e;
    ram_cell[     202] = 32'h0;  // 32'h9c5cc8d9;
    ram_cell[     203] = 32'h0;  // 32'h1b75fa4c;
    ram_cell[     204] = 32'h0;  // 32'h279be2f0;
    ram_cell[     205] = 32'h0;  // 32'hcee83a6f;
    ram_cell[     206] = 32'h0;  // 32'h20bc4c93;
    ram_cell[     207] = 32'h0;  // 32'ha5ef4d50;
    ram_cell[     208] = 32'h0;  // 32'h43a185bf;
    ram_cell[     209] = 32'h0;  // 32'hc260db92;
    ram_cell[     210] = 32'h0;  // 32'h8b5bca93;
    ram_cell[     211] = 32'h0;  // 32'h82fc729f;
    ram_cell[     212] = 32'h0;  // 32'h16a27b27;
    ram_cell[     213] = 32'h0;  // 32'h10d5344e;
    ram_cell[     214] = 32'h0;  // 32'h23b27124;
    ram_cell[     215] = 32'h0;  // 32'hb8cd229d;
    ram_cell[     216] = 32'h0;  // 32'he4457087;
    ram_cell[     217] = 32'h0;  // 32'h4f885d79;
    ram_cell[     218] = 32'h0;  // 32'h03195f47;
    ram_cell[     219] = 32'h0;  // 32'hdb3d2221;
    ram_cell[     220] = 32'h0;  // 32'h1acf9e0f;
    ram_cell[     221] = 32'h0;  // 32'h36cfb471;
    ram_cell[     222] = 32'h0;  // 32'h40d7d367;
    ram_cell[     223] = 32'h0;  // 32'h999de79e;
    ram_cell[     224] = 32'h0;  // 32'he1ebadb7;
    ram_cell[     225] = 32'h0;  // 32'h501c38e3;
    ram_cell[     226] = 32'h0;  // 32'h07c9251d;
    ram_cell[     227] = 32'h0;  // 32'hff72b949;
    ram_cell[     228] = 32'h0;  // 32'hdf24b5d5;
    ram_cell[     229] = 32'h0;  // 32'hec26ec45;
    ram_cell[     230] = 32'h0;  // 32'h82a305ec;
    ram_cell[     231] = 32'h0;  // 32'h67c95120;
    ram_cell[     232] = 32'h0;  // 32'h2e7ad8e7;
    ram_cell[     233] = 32'h0;  // 32'hacfea1a2;
    ram_cell[     234] = 32'h0;  // 32'h14e4b9b0;
    ram_cell[     235] = 32'h0;  // 32'he2c0f7ce;
    ram_cell[     236] = 32'h0;  // 32'h7b6a685b;
    ram_cell[     237] = 32'h0;  // 32'hc8f5301c;
    ram_cell[     238] = 32'h0;  // 32'h4a73ea7c;
    ram_cell[     239] = 32'h0;  // 32'h95a23f96;
    ram_cell[     240] = 32'h0;  // 32'hcbbb8a02;
    ram_cell[     241] = 32'h0;  // 32'h39f947d8;
    ram_cell[     242] = 32'h0;  // 32'h7eca0550;
    ram_cell[     243] = 32'h0;  // 32'hbd158ca7;
    ram_cell[     244] = 32'h0;  // 32'h59136c97;
    ram_cell[     245] = 32'h0;  // 32'h9e94fd7e;
    ram_cell[     246] = 32'h0;  // 32'h45877980;
    ram_cell[     247] = 32'h0;  // 32'h807225ac;
    ram_cell[     248] = 32'h0;  // 32'haaec9bbd;
    ram_cell[     249] = 32'h0;  // 32'hce1d667c;
    ram_cell[     250] = 32'h0;  // 32'hc2d78e25;
    ram_cell[     251] = 32'h0;  // 32'hb7c58eeb;
    ram_cell[     252] = 32'h0;  // 32'h1cd0c810;
    ram_cell[     253] = 32'h0;  // 32'h829f65ec;
    ram_cell[     254] = 32'h0;  // 32'h8c1b5d92;
    ram_cell[     255] = 32'h0;  // 32'he7e5ee8d;
    // src matrix A
    ram_cell[     256] = 32'hbc33052e;
    ram_cell[     257] = 32'h4a447e18;
    ram_cell[     258] = 32'h45e9e21f;
    ram_cell[     259] = 32'h4bb7a4e6;
    ram_cell[     260] = 32'ha98a0c51;
    ram_cell[     261] = 32'h8cafc001;
    ram_cell[     262] = 32'hbc5f0783;
    ram_cell[     263] = 32'h7887cd73;
    ram_cell[     264] = 32'h17ae6356;
    ram_cell[     265] = 32'hffb53f6f;
    ram_cell[     266] = 32'h7439a415;
    ram_cell[     267] = 32'h3c232384;
    ram_cell[     268] = 32'h3560b013;
    ram_cell[     269] = 32'hba327dda;
    ram_cell[     270] = 32'h9e1853b6;
    ram_cell[     271] = 32'h4749e3d2;
    ram_cell[     272] = 32'h47eaea72;
    ram_cell[     273] = 32'hb7fb33a0;
    ram_cell[     274] = 32'h31b0734c;
    ram_cell[     275] = 32'h0f6a4d63;
    ram_cell[     276] = 32'h5646d906;
    ram_cell[     277] = 32'hc14541f5;
    ram_cell[     278] = 32'h66f04dc2;
    ram_cell[     279] = 32'h27fb3db1;
    ram_cell[     280] = 32'hfc6338a5;
    ram_cell[     281] = 32'hca0e0582;
    ram_cell[     282] = 32'hcd4dc82c;
    ram_cell[     283] = 32'hbe3c1938;
    ram_cell[     284] = 32'h7a362577;
    ram_cell[     285] = 32'ha2597f9a;
    ram_cell[     286] = 32'hc84d597e;
    ram_cell[     287] = 32'he2099f27;
    ram_cell[     288] = 32'hbf7ac022;
    ram_cell[     289] = 32'he2f6a544;
    ram_cell[     290] = 32'h29745e13;
    ram_cell[     291] = 32'hafc16a1f;
    ram_cell[     292] = 32'h942159a0;
    ram_cell[     293] = 32'h4d092657;
    ram_cell[     294] = 32'hd7ba3c4a;
    ram_cell[     295] = 32'h31d5baf4;
    ram_cell[     296] = 32'hc0869ff4;
    ram_cell[     297] = 32'h31c31c52;
    ram_cell[     298] = 32'h397cbced;
    ram_cell[     299] = 32'h18620257;
    ram_cell[     300] = 32'hdc77ba25;
    ram_cell[     301] = 32'h8e5a30f7;
    ram_cell[     302] = 32'h46bbc120;
    ram_cell[     303] = 32'h60a2b08d;
    ram_cell[     304] = 32'h169330f9;
    ram_cell[     305] = 32'hc6947a0f;
    ram_cell[     306] = 32'h30844474;
    ram_cell[     307] = 32'h54ffa39e;
    ram_cell[     308] = 32'h4cd7e417;
    ram_cell[     309] = 32'h1f7b8d03;
    ram_cell[     310] = 32'h3bb0b7c1;
    ram_cell[     311] = 32'h00ba8e5d;
    ram_cell[     312] = 32'h6a52d2c8;
    ram_cell[     313] = 32'h84b814b0;
    ram_cell[     314] = 32'hb8ee1fd6;
    ram_cell[     315] = 32'h47380f43;
    ram_cell[     316] = 32'hb63b27da;
    ram_cell[     317] = 32'ha084e55c;
    ram_cell[     318] = 32'hb84d9f69;
    ram_cell[     319] = 32'hf1a86187;
    ram_cell[     320] = 32'h0e787638;
    ram_cell[     321] = 32'hdf4178c4;
    ram_cell[     322] = 32'h0e8bb539;
    ram_cell[     323] = 32'h6406e40f;
    ram_cell[     324] = 32'h2725da9b;
    ram_cell[     325] = 32'hfffb8d79;
    ram_cell[     326] = 32'h813fc90b;
    ram_cell[     327] = 32'hf4b0404a;
    ram_cell[     328] = 32'hfdbd18a7;
    ram_cell[     329] = 32'he7f2ded6;
    ram_cell[     330] = 32'ha82a8011;
    ram_cell[     331] = 32'h5eab04f3;
    ram_cell[     332] = 32'hf332a345;
    ram_cell[     333] = 32'h4ef47d8d;
    ram_cell[     334] = 32'hc0ca1b6a;
    ram_cell[     335] = 32'h7de59a20;
    ram_cell[     336] = 32'h7422b263;
    ram_cell[     337] = 32'h07cfe480;
    ram_cell[     338] = 32'haebd02e0;
    ram_cell[     339] = 32'hc52c0401;
    ram_cell[     340] = 32'ha9813c58;
    ram_cell[     341] = 32'h61ff2326;
    ram_cell[     342] = 32'h8d75b974;
    ram_cell[     343] = 32'h5170f14d;
    ram_cell[     344] = 32'hbc632f59;
    ram_cell[     345] = 32'he6e639df;
    ram_cell[     346] = 32'hd37f8f7e;
    ram_cell[     347] = 32'h124c9317;
    ram_cell[     348] = 32'h27792b59;
    ram_cell[     349] = 32'hc652ecfa;
    ram_cell[     350] = 32'hc5d5a7c5;
    ram_cell[     351] = 32'h8ce6bd02;
    ram_cell[     352] = 32'h61f54a65;
    ram_cell[     353] = 32'h1196ec2a;
    ram_cell[     354] = 32'h6ccca934;
    ram_cell[     355] = 32'h8a122c5d;
    ram_cell[     356] = 32'hef2728b1;
    ram_cell[     357] = 32'h0308f44d;
    ram_cell[     358] = 32'h0ad98303;
    ram_cell[     359] = 32'hee02a34b;
    ram_cell[     360] = 32'h6f49feb7;
    ram_cell[     361] = 32'h3ca775e3;
    ram_cell[     362] = 32'h6bf0169d;
    ram_cell[     363] = 32'hf9ee7ad7;
    ram_cell[     364] = 32'hca95b65f;
    ram_cell[     365] = 32'hc2912e4a;
    ram_cell[     366] = 32'ha4bec1ce;
    ram_cell[     367] = 32'h4ebf8de8;
    ram_cell[     368] = 32'h0a582b35;
    ram_cell[     369] = 32'h7d9ada54;
    ram_cell[     370] = 32'hf55a2813;
    ram_cell[     371] = 32'h1d946c34;
    ram_cell[     372] = 32'h0ab97f06;
    ram_cell[     373] = 32'hf2e1f7a5;
    ram_cell[     374] = 32'hecea06bc;
    ram_cell[     375] = 32'hf2e79515;
    ram_cell[     376] = 32'h80788981;
    ram_cell[     377] = 32'h0636abcb;
    ram_cell[     378] = 32'h324b4d88;
    ram_cell[     379] = 32'h928288a3;
    ram_cell[     380] = 32'h7081f5b4;
    ram_cell[     381] = 32'h4f74fc1b;
    ram_cell[     382] = 32'h6fa3f88b;
    ram_cell[     383] = 32'h98289dff;
    ram_cell[     384] = 32'h3b1abb4a;
    ram_cell[     385] = 32'h9d2c90a0;
    ram_cell[     386] = 32'h8b711faf;
    ram_cell[     387] = 32'h76927050;
    ram_cell[     388] = 32'h7fc70874;
    ram_cell[     389] = 32'h8fd35120;
    ram_cell[     390] = 32'h56ff3bcc;
    ram_cell[     391] = 32'h0a60ebfd;
    ram_cell[     392] = 32'h76378a3e;
    ram_cell[     393] = 32'h5da067d9;
    ram_cell[     394] = 32'h6f04b8fd;
    ram_cell[     395] = 32'h6f336c43;
    ram_cell[     396] = 32'he2d55f5b;
    ram_cell[     397] = 32'hae85e5c1;
    ram_cell[     398] = 32'h42d3b7c7;
    ram_cell[     399] = 32'h83509e7b;
    ram_cell[     400] = 32'hf6f1247a;
    ram_cell[     401] = 32'h2ff41261;
    ram_cell[     402] = 32'h6884dec3;
    ram_cell[     403] = 32'he2a9711c;
    ram_cell[     404] = 32'h56d8f79f;
    ram_cell[     405] = 32'h7cea3ee4;
    ram_cell[     406] = 32'h42db55ef;
    ram_cell[     407] = 32'he07621e1;
    ram_cell[     408] = 32'h1f682c68;
    ram_cell[     409] = 32'h80f865b2;
    ram_cell[     410] = 32'h791e227c;
    ram_cell[     411] = 32'h32a22e3f;
    ram_cell[     412] = 32'he7c081a5;
    ram_cell[     413] = 32'h19c00c20;
    ram_cell[     414] = 32'hbcedff70;
    ram_cell[     415] = 32'h9b65aa4b;
    ram_cell[     416] = 32'hd971fcd4;
    ram_cell[     417] = 32'hc558d2ba;
    ram_cell[     418] = 32'hed591a19;
    ram_cell[     419] = 32'h2bf80c0e;
    ram_cell[     420] = 32'h7abcb4b8;
    ram_cell[     421] = 32'h8fce27d4;
    ram_cell[     422] = 32'h2c2c6e6d;
    ram_cell[     423] = 32'h2b8b39d3;
    ram_cell[     424] = 32'h4789068d;
    ram_cell[     425] = 32'h4d2f82c5;
    ram_cell[     426] = 32'he7054238;
    ram_cell[     427] = 32'h586b996f;
    ram_cell[     428] = 32'h24babba2;
    ram_cell[     429] = 32'hc4e60f46;
    ram_cell[     430] = 32'h16e4815a;
    ram_cell[     431] = 32'h119eb823;
    ram_cell[     432] = 32'h12558af0;
    ram_cell[     433] = 32'h5da9ff16;
    ram_cell[     434] = 32'h97d5d9a8;
    ram_cell[     435] = 32'h3b24065a;
    ram_cell[     436] = 32'he4b2f904;
    ram_cell[     437] = 32'h318caacb;
    ram_cell[     438] = 32'h126ca504;
    ram_cell[     439] = 32'h2aa6a6d8;
    ram_cell[     440] = 32'h73a74681;
    ram_cell[     441] = 32'h6e03c132;
    ram_cell[     442] = 32'h69135a1d;
    ram_cell[     443] = 32'h16ebd155;
    ram_cell[     444] = 32'hddf56071;
    ram_cell[     445] = 32'h65e27f7f;
    ram_cell[     446] = 32'h63c3bda2;
    ram_cell[     447] = 32'h77f8b626;
    ram_cell[     448] = 32'h400cd41f;
    ram_cell[     449] = 32'h6a2576a3;
    ram_cell[     450] = 32'hdb79d163;
    ram_cell[     451] = 32'ha4eb8830;
    ram_cell[     452] = 32'hd51aa170;
    ram_cell[     453] = 32'hdcd3c473;
    ram_cell[     454] = 32'hca01204f;
    ram_cell[     455] = 32'hed18291f;
    ram_cell[     456] = 32'he3724afd;
    ram_cell[     457] = 32'he938a696;
    ram_cell[     458] = 32'hc43baa4a;
    ram_cell[     459] = 32'hdfc2d589;
    ram_cell[     460] = 32'h86ca62b2;
    ram_cell[     461] = 32'h6c0704b5;
    ram_cell[     462] = 32'hae01034b;
    ram_cell[     463] = 32'h59a54124;
    ram_cell[     464] = 32'h8f2ee969;
    ram_cell[     465] = 32'h9ca1542c;
    ram_cell[     466] = 32'hb479e2fd;
    ram_cell[     467] = 32'h377414da;
    ram_cell[     468] = 32'hec214638;
    ram_cell[     469] = 32'h56a22e58;
    ram_cell[     470] = 32'hded1059e;
    ram_cell[     471] = 32'hbfca2f59;
    ram_cell[     472] = 32'h10d5e9d1;
    ram_cell[     473] = 32'h6c67f461;
    ram_cell[     474] = 32'he3b2d4ae;
    ram_cell[     475] = 32'ha1020ccf;
    ram_cell[     476] = 32'h4859dd02;
    ram_cell[     477] = 32'hcb417f47;
    ram_cell[     478] = 32'h5ede9880;
    ram_cell[     479] = 32'hb7dfacde;
    ram_cell[     480] = 32'he0b5e906;
    ram_cell[     481] = 32'hf4b453eb;
    ram_cell[     482] = 32'h10118306;
    ram_cell[     483] = 32'h830b1c2b;
    ram_cell[     484] = 32'h452a10e5;
    ram_cell[     485] = 32'h8f25cf21;
    ram_cell[     486] = 32'h253ffd0b;
    ram_cell[     487] = 32'h8b9c363e;
    ram_cell[     488] = 32'h22f62ad2;
    ram_cell[     489] = 32'hcc2f3884;
    ram_cell[     490] = 32'hbcd0b4c9;
    ram_cell[     491] = 32'haa7c81f9;
    ram_cell[     492] = 32'hea00f209;
    ram_cell[     493] = 32'h2cdcfa43;
    ram_cell[     494] = 32'ha27410b0;
    ram_cell[     495] = 32'hd4ebee49;
    ram_cell[     496] = 32'h44065bf4;
    ram_cell[     497] = 32'hc5a4c70b;
    ram_cell[     498] = 32'ha746d203;
    ram_cell[     499] = 32'h56f7e84b;
    ram_cell[     500] = 32'h51c4e460;
    ram_cell[     501] = 32'h158861c6;
    ram_cell[     502] = 32'h07cd72ca;
    ram_cell[     503] = 32'h649f0592;
    ram_cell[     504] = 32'h5fcdca2f;
    ram_cell[     505] = 32'h85a8b09b;
    ram_cell[     506] = 32'h519badda;
    ram_cell[     507] = 32'h82d80614;
    ram_cell[     508] = 32'hca53cf7c;
    ram_cell[     509] = 32'hf20878ae;
    ram_cell[     510] = 32'hf1e7d6fa;
    ram_cell[     511] = 32'hb195052f;
    // src matrix B
    ram_cell[     512] = 32'hcb294291;
    ram_cell[     513] = 32'hfdc0845f;
    ram_cell[     514] = 32'hdcb47265;
    ram_cell[     515] = 32'h055803ce;
    ram_cell[     516] = 32'h7b0cd4e8;
    ram_cell[     517] = 32'h5811e17a;
    ram_cell[     518] = 32'h10f5d836;
    ram_cell[     519] = 32'hdaee8d77;
    ram_cell[     520] = 32'h83feb21f;
    ram_cell[     521] = 32'h1b6ce7fd;
    ram_cell[     522] = 32'hace653d1;
    ram_cell[     523] = 32'h944d4a05;
    ram_cell[     524] = 32'h97f79992;
    ram_cell[     525] = 32'h1e785b29;
    ram_cell[     526] = 32'hab1a4a6f;
    ram_cell[     527] = 32'hfa14f3a6;
    ram_cell[     528] = 32'h64d6fe85;
    ram_cell[     529] = 32'h7f9b75da;
    ram_cell[     530] = 32'h0b247b9c;
    ram_cell[     531] = 32'h897d59cd;
    ram_cell[     532] = 32'hc68da6d2;
    ram_cell[     533] = 32'he2e25ab2;
    ram_cell[     534] = 32'h85979337;
    ram_cell[     535] = 32'h522f03ed;
    ram_cell[     536] = 32'hc893c688;
    ram_cell[     537] = 32'h222772e1;
    ram_cell[     538] = 32'h490941a4;
    ram_cell[     539] = 32'hc21b6ac6;
    ram_cell[     540] = 32'hb031f8ca;
    ram_cell[     541] = 32'h1b23050b;
    ram_cell[     542] = 32'h83689bad;
    ram_cell[     543] = 32'hdf6afae6;
    ram_cell[     544] = 32'h66906109;
    ram_cell[     545] = 32'h7c4bc355;
    ram_cell[     546] = 32'h85d60c15;
    ram_cell[     547] = 32'h5728939e;
    ram_cell[     548] = 32'h2219ba09;
    ram_cell[     549] = 32'h26a4b793;
    ram_cell[     550] = 32'hd0c2192f;
    ram_cell[     551] = 32'hb26b4d00;
    ram_cell[     552] = 32'h131d89be;
    ram_cell[     553] = 32'h4e7e950f;
    ram_cell[     554] = 32'he0d4c165;
    ram_cell[     555] = 32'h2d220930;
    ram_cell[     556] = 32'h8f3b1378;
    ram_cell[     557] = 32'hba51cdaa;
    ram_cell[     558] = 32'h497eb6a1;
    ram_cell[     559] = 32'h24d7887d;
    ram_cell[     560] = 32'h152993b6;
    ram_cell[     561] = 32'h705ba580;
    ram_cell[     562] = 32'had15f9dd;
    ram_cell[     563] = 32'hbf43981d;
    ram_cell[     564] = 32'he53c083c;
    ram_cell[     565] = 32'hd608d242;
    ram_cell[     566] = 32'h0b395ddf;
    ram_cell[     567] = 32'he25deecf;
    ram_cell[     568] = 32'h0b69e45f;
    ram_cell[     569] = 32'h9be0c70b;
    ram_cell[     570] = 32'he3386184;
    ram_cell[     571] = 32'h237045cc;
    ram_cell[     572] = 32'h88ec8529;
    ram_cell[     573] = 32'h109c0dd0;
    ram_cell[     574] = 32'hfe8a38ae;
    ram_cell[     575] = 32'h92572943;
    ram_cell[     576] = 32'h994b8b62;
    ram_cell[     577] = 32'h280423f2;
    ram_cell[     578] = 32'h028f0faf;
    ram_cell[     579] = 32'h1ce3f3e7;
    ram_cell[     580] = 32'h270b7378;
    ram_cell[     581] = 32'h8cb8199e;
    ram_cell[     582] = 32'hed373f7b;
    ram_cell[     583] = 32'h8f21ce77;
    ram_cell[     584] = 32'h6c4fdabf;
    ram_cell[     585] = 32'h836949e6;
    ram_cell[     586] = 32'h4640f508;
    ram_cell[     587] = 32'h070bf071;
    ram_cell[     588] = 32'h6a23f5a8;
    ram_cell[     589] = 32'ha68f0bbb;
    ram_cell[     590] = 32'h01dbf550;
    ram_cell[     591] = 32'h31c9069f;
    ram_cell[     592] = 32'h8ae652fc;
    ram_cell[     593] = 32'hcc4ed57e;
    ram_cell[     594] = 32'ha39fb49f;
    ram_cell[     595] = 32'hbee7359f;
    ram_cell[     596] = 32'h7cf2f367;
    ram_cell[     597] = 32'hd4325798;
    ram_cell[     598] = 32'hf6928974;
    ram_cell[     599] = 32'h97e95d2d;
    ram_cell[     600] = 32'hf68c382e;
    ram_cell[     601] = 32'h7744d594;
    ram_cell[     602] = 32'h64554312;
    ram_cell[     603] = 32'h0e27b18f;
    ram_cell[     604] = 32'hbe04a233;
    ram_cell[     605] = 32'h4cb9f9b5;
    ram_cell[     606] = 32'h61864c9c;
    ram_cell[     607] = 32'hb09fa490;
    ram_cell[     608] = 32'hf244dddd;
    ram_cell[     609] = 32'ha530b271;
    ram_cell[     610] = 32'h17976ef3;
    ram_cell[     611] = 32'h667b6bcf;
    ram_cell[     612] = 32'h0621a4ad;
    ram_cell[     613] = 32'h354327b6;
    ram_cell[     614] = 32'h76d50e15;
    ram_cell[     615] = 32'h31134b5e;
    ram_cell[     616] = 32'hbb862091;
    ram_cell[     617] = 32'h501e2093;
    ram_cell[     618] = 32'he3186a23;
    ram_cell[     619] = 32'hb3883f4e;
    ram_cell[     620] = 32'h0509f8c7;
    ram_cell[     621] = 32'h8849ea89;
    ram_cell[     622] = 32'hf55cfc5c;
    ram_cell[     623] = 32'h4e1ca36f;
    ram_cell[     624] = 32'h8fd8179b;
    ram_cell[     625] = 32'h0f9925ec;
    ram_cell[     626] = 32'h97e1293c;
    ram_cell[     627] = 32'h0a9f990a;
    ram_cell[     628] = 32'ha395b265;
    ram_cell[     629] = 32'h8639aebf;
    ram_cell[     630] = 32'h789f33e9;
    ram_cell[     631] = 32'h42dbc8e8;
    ram_cell[     632] = 32'h6374287e;
    ram_cell[     633] = 32'h9ede355c;
    ram_cell[     634] = 32'hebddb007;
    ram_cell[     635] = 32'h1461d708;
    ram_cell[     636] = 32'he2a846f9;
    ram_cell[     637] = 32'h93c3449c;
    ram_cell[     638] = 32'hcb520089;
    ram_cell[     639] = 32'hb58b15f4;
    ram_cell[     640] = 32'h713b16d3;
    ram_cell[     641] = 32'h510bf733;
    ram_cell[     642] = 32'h3c6b1ddb;
    ram_cell[     643] = 32'h1f12ca13;
    ram_cell[     644] = 32'h73e4ebde;
    ram_cell[     645] = 32'h7fd5ffd8;
    ram_cell[     646] = 32'h69f9c9b4;
    ram_cell[     647] = 32'h1c94c47a;
    ram_cell[     648] = 32'h09634ae6;
    ram_cell[     649] = 32'he7d58bdd;
    ram_cell[     650] = 32'h6940186a;
    ram_cell[     651] = 32'h42986e83;
    ram_cell[     652] = 32'h079e6e32;
    ram_cell[     653] = 32'hd2751d02;
    ram_cell[     654] = 32'h48a097ae;
    ram_cell[     655] = 32'h218e725b;
    ram_cell[     656] = 32'h1bad3a77;
    ram_cell[     657] = 32'h2f314ebc;
    ram_cell[     658] = 32'h1ad8d3d0;
    ram_cell[     659] = 32'h800a330b;
    ram_cell[     660] = 32'hb839ecb2;
    ram_cell[     661] = 32'hacde5351;
    ram_cell[     662] = 32'hf60d0487;
    ram_cell[     663] = 32'h92036948;
    ram_cell[     664] = 32'h97a36ba3;
    ram_cell[     665] = 32'h1c79f2ce;
    ram_cell[     666] = 32'h1a01b26d;
    ram_cell[     667] = 32'h51d738f2;
    ram_cell[     668] = 32'h086139ce;
    ram_cell[     669] = 32'he0466f26;
    ram_cell[     670] = 32'h8daad142;
    ram_cell[     671] = 32'hc37a747a;
    ram_cell[     672] = 32'hc1a8f0b1;
    ram_cell[     673] = 32'hd2155f07;
    ram_cell[     674] = 32'h10223839;
    ram_cell[     675] = 32'h50c149f3;
    ram_cell[     676] = 32'h3d48ad54;
    ram_cell[     677] = 32'h7f01aaf6;
    ram_cell[     678] = 32'hb62cac92;
    ram_cell[     679] = 32'h56c0b22f;
    ram_cell[     680] = 32'h73dd2304;
    ram_cell[     681] = 32'hb6e589d4;
    ram_cell[     682] = 32'h0b6e333a;
    ram_cell[     683] = 32'he1325237;
    ram_cell[     684] = 32'h976949d6;
    ram_cell[     685] = 32'h0497cdbc;
    ram_cell[     686] = 32'hd26ea500;
    ram_cell[     687] = 32'hb3b6719b;
    ram_cell[     688] = 32'h8b5ca312;
    ram_cell[     689] = 32'he7e1e0c0;
    ram_cell[     690] = 32'hf09b4646;
    ram_cell[     691] = 32'h055c3350;
    ram_cell[     692] = 32'h4ab51172;
    ram_cell[     693] = 32'hde898cc1;
    ram_cell[     694] = 32'he0343605;
    ram_cell[     695] = 32'h66dd91ff;
    ram_cell[     696] = 32'h68443087;
    ram_cell[     697] = 32'h06025005;
    ram_cell[     698] = 32'hf87a64aa;
    ram_cell[     699] = 32'hf9b14d57;
    ram_cell[     700] = 32'h95a47cc1;
    ram_cell[     701] = 32'h78cd0a82;
    ram_cell[     702] = 32'hc255f4ee;
    ram_cell[     703] = 32'h800d7e1e;
    ram_cell[     704] = 32'hfb2152e4;
    ram_cell[     705] = 32'h269e8d70;
    ram_cell[     706] = 32'h20989a1f;
    ram_cell[     707] = 32'h3bbb2373;
    ram_cell[     708] = 32'h2b407996;
    ram_cell[     709] = 32'h7eaa30ce;
    ram_cell[     710] = 32'hd7a23833;
    ram_cell[     711] = 32'h40a3c19d;
    ram_cell[     712] = 32'hed1a51a8;
    ram_cell[     713] = 32'h4de7b8bd;
    ram_cell[     714] = 32'hb9d2526f;
    ram_cell[     715] = 32'h2f26245e;
    ram_cell[     716] = 32'h8bc30cd7;
    ram_cell[     717] = 32'h64a25607;
    ram_cell[     718] = 32'hd80e3d05;
    ram_cell[     719] = 32'h689284a8;
    ram_cell[     720] = 32'hf6f27a82;
    ram_cell[     721] = 32'h8dee611f;
    ram_cell[     722] = 32'h12d3aada;
    ram_cell[     723] = 32'hdbdebff7;
    ram_cell[     724] = 32'hd183323f;
    ram_cell[     725] = 32'h88edb21c;
    ram_cell[     726] = 32'h60b5c35e;
    ram_cell[     727] = 32'hefedd23d;
    ram_cell[     728] = 32'h021a55d0;
    ram_cell[     729] = 32'h9afd1aaf;
    ram_cell[     730] = 32'h55cc612f;
    ram_cell[     731] = 32'he56472d0;
    ram_cell[     732] = 32'h4be43ffd;
    ram_cell[     733] = 32'ha1b8b0b4;
    ram_cell[     734] = 32'hba5cf3f8;
    ram_cell[     735] = 32'he853c380;
    ram_cell[     736] = 32'h07641f49;
    ram_cell[     737] = 32'h09bb6ccb;
    ram_cell[     738] = 32'h412ea5b9;
    ram_cell[     739] = 32'h2d1d830a;
    ram_cell[     740] = 32'h587f8d36;
    ram_cell[     741] = 32'hf3332bcf;
    ram_cell[     742] = 32'h5e357c39;
    ram_cell[     743] = 32'ha4a11319;
    ram_cell[     744] = 32'h6fc8603a;
    ram_cell[     745] = 32'hc4228a85;
    ram_cell[     746] = 32'haa6eda42;
    ram_cell[     747] = 32'hc21e91b4;
    ram_cell[     748] = 32'h56331d5d;
    ram_cell[     749] = 32'h74ad6a53;
    ram_cell[     750] = 32'h3a112fa3;
    ram_cell[     751] = 32'hff62a8a3;
    ram_cell[     752] = 32'h62e09c1c;
    ram_cell[     753] = 32'hc3a4a70e;
    ram_cell[     754] = 32'he1d0d30d;
    ram_cell[     755] = 32'h4de3348d;
    ram_cell[     756] = 32'hac3b341a;
    ram_cell[     757] = 32'h99304536;
    ram_cell[     758] = 32'hf49197b4;
    ram_cell[     759] = 32'h5b682516;
    ram_cell[     760] = 32'h2405258d;
    ram_cell[     761] = 32'he90749be;
    ram_cell[     762] = 32'hb653a0a5;
    ram_cell[     763] = 32'h10536de6;
    ram_cell[     764] = 32'hebb749b3;
    ram_cell[     765] = 32'hacc1ecad;
    ram_cell[     766] = 32'h6c21530c;
    ram_cell[     767] = 32'h35a8956c;
end

endmodule

