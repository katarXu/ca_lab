
module mem #(                   // 
    parameter  ADDR_LEN  = 11   // 
) (
    input  clk, rst,
    input  [ADDR_LEN-1:0] addr, // memory address
    output reg [31:0] rd_data,  // data read out
    input  wr_req,
    input  [31:0] wr_data       // data write in
);
localparam MEM_SIZE = 1<<ADDR_LEN;
reg [31:0] ram_cell [2000];

always @ (posedge clk or posedge rst)
    if(rst)
        rd_data <= 0;
    else
        rd_data <= ram_cell[addr];

always @ (posedge clk)
    if(wr_req) 
        ram_cell[addr] <= wr_data;

initial begin
    /*
    ram_cell[       0] = 32'h0000005e;
    ram_cell[       1] = 32'h000000b8;
    ram_cell[       2] = 32'h00000051;
    ram_cell[       3] = 32'h00000021;
    ram_cell[       4] = 32'h000000ff;
    ram_cell[       5] = 32'h0000007a;
    ram_cell[       6] = 32'h00000033;
    ram_cell[       7] = 32'h000000e4;
    ram_cell[       8] = 32'h000000fa;
    ram_cell[       9] = 32'h0000004e;
    ram_cell[      10] = 32'h000000c0;
    ram_cell[      11] = 32'h00000093;
    ram_cell[      12] = 32'h000000bb;
    ram_cell[      13] = 32'h000000e9;
    ram_cell[      14] = 32'h00000041;
    ram_cell[      15] = 32'h00000081;
    ram_cell[      16] = 32'h0000007f;
    ram_cell[      17] = 32'h000000c5;
    ram_cell[      18] = 32'h000000f6;
    ram_cell[      19] = 32'h000000bc;
    ram_cell[      20] = 32'h00000012;
    ram_cell[      21] = 32'h000000a0;
    ram_cell[      22] = 32'h00000001;
    ram_cell[      23] = 32'h0000009d;
    ram_cell[      24] = 32'h000000e7;
    ram_cell[      25] = 32'h0000000b;
    ram_cell[      26] = 32'h000000cb;
    ram_cell[      27] = 32'h000000cd;
    ram_cell[      28] = 32'h000000cf;
    ram_cell[      29] = 32'h00000044;
    ram_cell[      30] = 32'h000000cc;
    ram_cell[      31] = 32'h000000ef;
    ram_cell[      32] = 32'h00000056;
    ram_cell[      33] = 32'h00000049;
    ram_cell[      34] = 32'h00000064;
    ram_cell[      35] = 32'h0000006e;
    ram_cell[      36] = 32'h0000003a;
    ram_cell[      37] = 32'h000000ed;
    ram_cell[      38] = 32'h00000009;
    ram_cell[      39] = 32'h000000f4;
    ram_cell[      40] = 32'h000000ec;
    ram_cell[      41] = 32'h0000005c;
    ram_cell[      42] = 32'h000000e1;
    ram_cell[      43] = 32'h00000032;
    ram_cell[      44] = 32'h000000ba;
    ram_cell[      45] = 32'h00000077;
    ram_cell[      46] = 32'h000000fb;
    ram_cell[      47] = 32'h000000e5;
    ram_cell[      48] = 32'h00000070;
    ram_cell[      49] = 32'h00000019;
    ram_cell[      50] = 32'h0000000a;
    ram_cell[      51] = 32'h00000010;
    ram_cell[      52] = 32'h000000d6;
    ram_cell[      53] = 32'h000000b6;
    ram_cell[      54] = 32'h000000a7;
    ram_cell[      55] = 32'h000000d1;
    ram_cell[      56] = 32'h0000003e;
    ram_cell[      57] = 32'h0000007b;
    ram_cell[      58] = 32'h0000006f;
    ram_cell[      59] = 32'h0000006b;
    ram_cell[      60] = 32'h00000060;
    ram_cell[      61] = 32'h000000f9;
    ram_cell[      62] = 32'h000000c7;
    ram_cell[      63] = 32'h00000075;
    ram_cell[      64] = 32'h00000066;
    ram_cell[      65] = 32'h0000004b;
    ram_cell[      66] = 32'h00000072;
    ram_cell[      67] = 32'h0000001f;
    ram_cell[      68] = 32'h00000050;
    ram_cell[      69] = 32'h00000038;
    ram_cell[      70] = 32'h00000020;
    ram_cell[      71] = 32'h00000025;
    ram_cell[      72] = 32'h00000024;
    ram_cell[      73] = 32'h00000018;
    ram_cell[      74] = 32'h00000095;
    ram_cell[      75] = 32'h000000f1;
    ram_cell[      76] = 32'h00000026;
    ram_cell[      77] = 32'h00000062;
    ram_cell[      78] = 32'h00000089;
    ram_cell[      79] = 32'h0000003d;
    ram_cell[      80] = 32'h00000014;
    ram_cell[      81] = 32'h00000039;
    ram_cell[      82] = 32'h000000be;
    ram_cell[      83] = 32'h0000002c;
    ram_cell[      84] = 32'h000000ca;
    ram_cell[      85] = 32'h0000008a;
    ram_cell[      86] = 32'h000000a8;
    ram_cell[      87] = 32'h000000e2;
    ram_cell[      88] = 32'h000000f3;
    ram_cell[      89] = 32'h00000022;
    ram_cell[      90] = 32'h000000de;
    ram_cell[      91] = 32'h00000091;
    ram_cell[      92] = 32'h00000076;
    ram_cell[      93] = 32'h000000e0;
    ram_cell[      94] = 32'h00000073;
    ram_cell[      95] = 32'h00000085;
    ram_cell[      96] = 32'h000000e6;
    ram_cell[      97] = 32'h000000eb;
    ram_cell[      98] = 32'h00000040;
    ram_cell[      99] = 32'h000000fe;
    ram_cell[     100] = 32'h00000046;
    ram_cell[     101] = 32'h00000058;
    ram_cell[     102] = 32'h000000af;
    ram_cell[     103] = 32'h00000068;
    ram_cell[     104] = 32'h00000084;
    ram_cell[     105] = 32'h00000088;
    ram_cell[     106] = 32'h00000047;
    ram_cell[     107] = 32'h000000b5;
    ram_cell[     108] = 32'h00000029;
    ram_cell[     109] = 32'h00000074;
    ram_cell[     110] = 32'h00000005;
    ram_cell[     111] = 32'h000000a1;
    ram_cell[     112] = 32'h0000008c;
    ram_cell[     113] = 32'h00000099;
    ram_cell[     114] = 32'h000000b3;
    ram_cell[     115] = 32'h000000f5;
    ram_cell[     116] = 32'h00000092;
    ram_cell[     117] = 32'h000000b4;
    ram_cell[     118] = 32'h0000001b;
    ram_cell[     119] = 32'h000000d3;
    ram_cell[     120] = 32'h000000fc;
    ram_cell[     121] = 32'h000000f0;
    ram_cell[     122] = 32'h00000006;
    ram_cell[     123] = 32'h000000ad;
    ram_cell[     124] = 32'h000000a5;
    ram_cell[     125] = 32'h000000aa;
    ram_cell[     126] = 32'h00000003;
    ram_cell[     127] = 32'h00000061;
    ram_cell[     128] = 32'h0000005d;
    ram_cell[     129] = 32'h000000d2;
    ram_cell[     130] = 32'h00000082;
    ram_cell[     131] = 32'h00000055;
    ram_cell[     132] = 32'h00000002;
    ram_cell[     133] = 32'h0000005f;
    ram_cell[     134] = 32'h0000003b;
    ram_cell[     135] = 32'h00000017;
    ram_cell[     136] = 32'h00000067;
    ram_cell[     137] = 32'h0000004c;
    ram_cell[     138] = 32'h0000001d;
    ram_cell[     139] = 32'h000000c8;
    ram_cell[     140] = 32'h000000dd;
    ram_cell[     141] = 32'h000000db;
    ram_cell[     142] = 32'h000000d0;
    ram_cell[     143] = 32'h0000009a;
    ram_cell[     144] = 32'h00000079;
    ram_cell[     145] = 32'h000000f2;
    ram_cell[     146] = 32'h00000057;
    ram_cell[     147] = 32'h00000035;
    ram_cell[     148] = 32'h0000004f;
    ram_cell[     149] = 32'h000000df;
    ram_cell[     150] = 32'h00000097;
    ram_cell[     151] = 32'h0000007c;
    ram_cell[     152] = 32'h0000005a;
    ram_cell[     153] = 32'h0000002d;
    ram_cell[     154] = 32'h000000a9;
    ram_cell[     155] = 32'h00000071;
    ram_cell[     156] = 32'h0000009f;
    ram_cell[     157] = 32'h00000090;
    ram_cell[     158] = 32'h000000bd;
    ram_cell[     159] = 32'h000000a4;
    ram_cell[     160] = 32'h0000002e;
    ram_cell[     161] = 32'h0000008e;
    ram_cell[     162] = 32'h0000008d;
    ram_cell[     163] = 32'h00000054;
    ram_cell[     164] = 32'h0000009b;
    ram_cell[     165] = 32'h00000043;
    ram_cell[     166] = 32'h00000094;
    ram_cell[     167] = 32'h000000f8;
    ram_cell[     168] = 32'h00000087;
    ram_cell[     169] = 32'h0000004d;
    ram_cell[     170] = 32'h0000000d;
    ram_cell[     171] = 32'h00000013;
    ram_cell[     172] = 32'h000000da;
    ram_cell[     173] = 32'h0000003f;
    ram_cell[     174] = 32'h0000007e;
    ram_cell[     175] = 32'h000000ac;
    ram_cell[     176] = 32'h000000e8;
    ram_cell[     177] = 32'h0000006c;
    ram_cell[     178] = 32'h00000083;
    ram_cell[     179] = 32'h000000b1;
    ram_cell[     180] = 32'h000000b7;
    ram_cell[     181] = 32'h000000bf;
    ram_cell[     182] = 32'h000000ea;
    ram_cell[     183] = 32'h00000078;
    ram_cell[     184] = 32'h00000027;
    ram_cell[     185] = 32'h0000002a;
    ram_cell[     186] = 32'h0000001a;
    ram_cell[     187] = 32'h000000a3;
    ram_cell[     188] = 32'h0000002f;
    ram_cell[     189] = 32'h000000c6;
    ram_cell[     190] = 32'h00000053;
    ram_cell[     191] = 32'h000000d9;
    ram_cell[     192] = 32'h000000b9;
    ram_cell[     193] = 32'h00000030;
    ram_cell[     194] = 32'h0000001c;
    ram_cell[     195] = 32'h00000028;
    ram_cell[     196] = 32'h00000037;
    ram_cell[     197] = 32'h000000b2;
    ram_cell[     198] = 32'h0000006d;
    ram_cell[     199] = 32'h00000036;
    ram_cell[     200] = 32'h000000e3;
    ram_cell[     201] = 32'h000000d7;
    ram_cell[     202] = 32'h00000096;
    ram_cell[     203] = 32'h000000c1;
    ram_cell[     204] = 32'h0000006a;
    ram_cell[     205] = 32'h00000016;
    ram_cell[     206] = 32'h0000008b;
    ram_cell[     207] = 32'h00000063;
    ram_cell[     208] = 32'h00000031;
    ram_cell[     209] = 32'h000000dc;
    ram_cell[     210] = 32'h000000ae;
    ram_cell[     211] = 32'h000000c2;
    ram_cell[     212] = 32'h000000c9;
    ram_cell[     213] = 32'h0000008f;
    ram_cell[     214] = 32'h000000a2;
    ram_cell[     215] = 32'h000000a6;
    ram_cell[     216] = 32'h00000065;
    ram_cell[     217] = 32'h000000c3;
    ram_cell[     218] = 32'h000000ee;
    ram_cell[     219] = 32'h0000000c;
    ram_cell[     220] = 32'h00000098;
    ram_cell[     221] = 32'h00000034;
    ram_cell[     222] = 32'h000000d5;
    ram_cell[     223] = 32'h00000004;
    ram_cell[     224] = 32'h0000005b;
    ram_cell[     225] = 32'h00000011;
    ram_cell[     226] = 32'h000000ce;
    ram_cell[     227] = 32'h00000000;
    ram_cell[     228] = 32'h0000001e;
    ram_cell[     229] = 32'h0000004a;
    ram_cell[     230] = 32'h0000003c;
    ram_cell[     231] = 32'h000000f7;
    ram_cell[     232] = 32'h000000c4;
    ram_cell[     233] = 32'h0000007d;
    ram_cell[     234] = 32'h00000048;
    ram_cell[     235] = 32'h000000d4;
    ram_cell[     236] = 32'h00000069;
    ram_cell[     237] = 32'h00000007;
    ram_cell[     238] = 32'h00000080;
    ram_cell[     239] = 32'h0000000f;
    ram_cell[     240] = 32'h00000045;
    ram_cell[     241] = 32'h0000000e;
    ram_cell[     242] = 32'h0000002b;
    ram_cell[     243] = 32'h000000ab;
    ram_cell[     244] = 32'h0000009e;
    ram_cell[     245] = 32'h000000b0;
    ram_cell[     246] = 32'h00000042;
    ram_cell[     247] = 32'h00000015;
    ram_cell[     248] = 32'h00000052;
    ram_cell[     249] = 32'h00000008;
    ram_cell[     250] = 32'h00000023;
    ram_cell[     251] = 32'h000000fd;
    ram_cell[     252] = 32'h00000059;
    ram_cell[     253] = 32'h0000009c;
    ram_cell[     254] = 32'h00000086;
    ram_cell[     255] = 32'h000000d8;
    */

    // dst matrix C
    ram_cell[       0] = 32'h0;  // 32'hc8528b48;
    ram_cell[       1] = 32'h0;  // 32'h45fe0cc5;
    ram_cell[       2] = 32'h0;  // 32'h437d9d40;
    ram_cell[       3] = 32'h0;  // 32'h394fa298;
    ram_cell[       4] = 32'h0;  // 32'hf296448e;
    ram_cell[       5] = 32'h0;  // 32'h9d60cdfb;
    ram_cell[       6] = 32'h0;  // 32'h64d460f0;
    ram_cell[       7] = 32'h0;  // 32'h9aeb3e36;
    ram_cell[       8] = 32'h0;  // 32'hcd02889d;
    ram_cell[       9] = 32'h0;  // 32'h951f7399;
    ram_cell[      10] = 32'h0;  // 32'h687eee57;
    ram_cell[      11] = 32'h0;  // 32'hc206a10e;
    ram_cell[      12] = 32'h0;  // 32'hbeecc07d;
    ram_cell[      13] = 32'h0;  // 32'h6c2754fb;
    ram_cell[      14] = 32'h0;  // 32'hff4f1b63;
    ram_cell[      15] = 32'h0;  // 32'h6a5f3004;
    ram_cell[      16] = 32'h0;  // 32'h497979cc;
    ram_cell[      17] = 32'h0;  // 32'hfae48e40;
    ram_cell[      18] = 32'h0;  // 32'h18ca6b5d;
    ram_cell[      19] = 32'h0;  // 32'h0723e7a1;
    ram_cell[      20] = 32'h0;  // 32'h3a0b46f4;
    ram_cell[      21] = 32'h0;  // 32'hf286bd18;
    ram_cell[      22] = 32'h0;  // 32'he1981f2f;
    ram_cell[      23] = 32'h0;  // 32'h84c0ad50;
    ram_cell[      24] = 32'h0;  // 32'hfab9802d;
    ram_cell[      25] = 32'h0;  // 32'h1ff1a4a5;
    ram_cell[      26] = 32'h0;  // 32'h3002e0af;
    ram_cell[      27] = 32'h0;  // 32'h80e90dd1;
    ram_cell[      28] = 32'h0;  // 32'hf42c91bd;
    ram_cell[      29] = 32'h0;  // 32'h64be79bc;
    ram_cell[      30] = 32'h0;  // 32'h854a3b0e;
    ram_cell[      31] = 32'h0;  // 32'h272c0da7;
    ram_cell[      32] = 32'h0;  // 32'h256a72d5;
    ram_cell[      33] = 32'h0;  // 32'hba49069a;
    ram_cell[      34] = 32'h0;  // 32'hce6f6b20;
    ram_cell[      35] = 32'h0;  // 32'h31cc0112;
    ram_cell[      36] = 32'h0;  // 32'hfd838b4c;
    ram_cell[      37] = 32'h0;  // 32'h3baceabb;
    ram_cell[      38] = 32'h0;  // 32'hccc3f923;
    ram_cell[      39] = 32'h0;  // 32'h307832fa;
    ram_cell[      40] = 32'h0;  // 32'h7cfbf780;
    ram_cell[      41] = 32'h0;  // 32'h4deef87c;
    ram_cell[      42] = 32'h0;  // 32'hc1f36df7;
    ram_cell[      43] = 32'h0;  // 32'h636e150b;
    ram_cell[      44] = 32'h0;  // 32'he4e3c00d;
    ram_cell[      45] = 32'h0;  // 32'h86ef543a;
    ram_cell[      46] = 32'h0;  // 32'hebf56b31;
    ram_cell[      47] = 32'h0;  // 32'h68095b4b;
    ram_cell[      48] = 32'h0;  // 32'h0995a617;
    ram_cell[      49] = 32'h0;  // 32'hed924fc7;
    ram_cell[      50] = 32'h0;  // 32'hd1ef9768;
    ram_cell[      51] = 32'h0;  // 32'h8df02f49;
    ram_cell[      52] = 32'h0;  // 32'h99763233;
    ram_cell[      53] = 32'h0;  // 32'h611b6901;
    ram_cell[      54] = 32'h0;  // 32'h05716fa1;
    ram_cell[      55] = 32'h0;  // 32'h3b4f9ee3;
    ram_cell[      56] = 32'h0;  // 32'h0bb4f1bb;
    ram_cell[      57] = 32'h0;  // 32'h2ac343aa;
    ram_cell[      58] = 32'h0;  // 32'h374d4816;
    ram_cell[      59] = 32'h0;  // 32'haf6c48e7;
    ram_cell[      60] = 32'h0;  // 32'h92f192ac;
    ram_cell[      61] = 32'h0;  // 32'haed715f2;
    ram_cell[      62] = 32'h0;  // 32'heff714be;
    ram_cell[      63] = 32'h0;  // 32'h9f4b9f45;
    ram_cell[      64] = 32'h0;  // 32'h9cadfad6;
    ram_cell[      65] = 32'h0;  // 32'h5a6101ee;
    ram_cell[      66] = 32'h0;  // 32'h5cdf0d9b;
    ram_cell[      67] = 32'h0;  // 32'hb710fc53;
    ram_cell[      68] = 32'h0;  // 32'hbc49b1d0;
    ram_cell[      69] = 32'h0;  // 32'h7f07b23a;
    ram_cell[      70] = 32'h0;  // 32'h2a772e1e;
    ram_cell[      71] = 32'h0;  // 32'h4f711a51;
    ram_cell[      72] = 32'h0;  // 32'h08d963e5;
    ram_cell[      73] = 32'h0;  // 32'h90d0c73b;
    ram_cell[      74] = 32'h0;  // 32'h757a54db;
    ram_cell[      75] = 32'h0;  // 32'h2970b4a7;
    ram_cell[      76] = 32'h0;  // 32'he2a71ada;
    ram_cell[      77] = 32'h0;  // 32'h4cd517c8;
    ram_cell[      78] = 32'h0;  // 32'h4701a18e;
    ram_cell[      79] = 32'h0;  // 32'h1c57a484;
    ram_cell[      80] = 32'h0;  // 32'h6ef874e2;
    ram_cell[      81] = 32'h0;  // 32'h14ffa445;
    ram_cell[      82] = 32'h0;  // 32'h2a54f25d;
    ram_cell[      83] = 32'h0;  // 32'h5039fe91;
    ram_cell[      84] = 32'h0;  // 32'he4812edd;
    ram_cell[      85] = 32'h0;  // 32'hc5ebf26f;
    ram_cell[      86] = 32'h0;  // 32'ha81394c3;
    ram_cell[      87] = 32'h0;  // 32'h195d47af;
    ram_cell[      88] = 32'h0;  // 32'h1d570290;
    ram_cell[      89] = 32'h0;  // 32'h5613aa8b;
    ram_cell[      90] = 32'h0;  // 32'h72278baf;
    ram_cell[      91] = 32'h0;  // 32'hb07009cb;
    ram_cell[      92] = 32'h0;  // 32'h5ac498e9;
    ram_cell[      93] = 32'h0;  // 32'h8d6de47d;
    ram_cell[      94] = 32'h0;  // 32'h724618ad;
    ram_cell[      95] = 32'h0;  // 32'h3187d9d3;
    ram_cell[      96] = 32'h0;  // 32'ha30c2d95;
    ram_cell[      97] = 32'h0;  // 32'hadbd93e7;
    ram_cell[      98] = 32'h0;  // 32'he6a2a278;
    ram_cell[      99] = 32'h0;  // 32'hb6c8055a;
    ram_cell[     100] = 32'h0;  // 32'h7f65c1cd;
    ram_cell[     101] = 32'h0;  // 32'hf86f21ff;
    ram_cell[     102] = 32'h0;  // 32'h63ff3be3;
    ram_cell[     103] = 32'h0;  // 32'hc098fce3;
    ram_cell[     104] = 32'h0;  // 32'h45a14b39;
    ram_cell[     105] = 32'h0;  // 32'h847b468b;
    ram_cell[     106] = 32'h0;  // 32'h2eeeecd4;
    ram_cell[     107] = 32'h0;  // 32'h63504c2e;
    ram_cell[     108] = 32'h0;  // 32'h89cb2d90;
    ram_cell[     109] = 32'h0;  // 32'hab2c26fc;
    ram_cell[     110] = 32'h0;  // 32'h516312c8;
    ram_cell[     111] = 32'h0;  // 32'hd89f0123;
    ram_cell[     112] = 32'h0;  // 32'hfdf06534;
    ram_cell[     113] = 32'h0;  // 32'h91c012b2;
    ram_cell[     114] = 32'h0;  // 32'hdfee8bf2;
    ram_cell[     115] = 32'h0;  // 32'h8d3fa35d;
    ram_cell[     116] = 32'h0;  // 32'h224d7e9b;
    ram_cell[     117] = 32'h0;  // 32'hfb3eb61c;
    ram_cell[     118] = 32'h0;  // 32'h5130abe6;
    ram_cell[     119] = 32'h0;  // 32'h5e5a6435;
    ram_cell[     120] = 32'h0;  // 32'hde3e36a9;
    ram_cell[     121] = 32'h0;  // 32'h5abcb5e0;
    ram_cell[     122] = 32'h0;  // 32'h0e855b85;
    ram_cell[     123] = 32'h0;  // 32'h1cd28488;
    ram_cell[     124] = 32'h0;  // 32'h7ba74598;
    ram_cell[     125] = 32'h0;  // 32'hb60df937;
    ram_cell[     126] = 32'h0;  // 32'hc41c78c3;
    ram_cell[     127] = 32'h0;  // 32'h47d28517;
    ram_cell[     128] = 32'h0;  // 32'h38ec48ca;
    ram_cell[     129] = 32'h0;  // 32'h849eff7a;
    ram_cell[     130] = 32'h0;  // 32'hb1ef4794;
    ram_cell[     131] = 32'h0;  // 32'h3a57b534;
    ram_cell[     132] = 32'h0;  // 32'h6e11364d;
    ram_cell[     133] = 32'h0;  // 32'ha74f25e6;
    ram_cell[     134] = 32'h0;  // 32'hf38aa065;
    ram_cell[     135] = 32'h0;  // 32'hf84b7b9b;
    ram_cell[     136] = 32'h0;  // 32'h1fe03dae;
    ram_cell[     137] = 32'h0;  // 32'had3d0143;
    ram_cell[     138] = 32'h0;  // 32'h9b6db6e0;
    ram_cell[     139] = 32'h0;  // 32'hd97b6b8f;
    ram_cell[     140] = 32'h0;  // 32'hd3775338;
    ram_cell[     141] = 32'h0;  // 32'h8eb52273;
    ram_cell[     142] = 32'h0;  // 32'h4e0b3d53;
    ram_cell[     143] = 32'h0;  // 32'hbcb19c47;
    ram_cell[     144] = 32'h0;  // 32'h073b05ea;
    ram_cell[     145] = 32'h0;  // 32'h3ce93c25;
    ram_cell[     146] = 32'h0;  // 32'h0987e271;
    ram_cell[     147] = 32'h0;  // 32'ha24ba13c;
    ram_cell[     148] = 32'h0;  // 32'h5ae19d12;
    ram_cell[     149] = 32'h0;  // 32'ha82c8dc5;
    ram_cell[     150] = 32'h0;  // 32'h2faaf83c;
    ram_cell[     151] = 32'h0;  // 32'hac197119;
    ram_cell[     152] = 32'h0;  // 32'ha145911a;
    ram_cell[     153] = 32'h0;  // 32'h810e665c;
    ram_cell[     154] = 32'h0;  // 32'h4d1a8dd5;
    ram_cell[     155] = 32'h0;  // 32'h622057e6;
    ram_cell[     156] = 32'h0;  // 32'h462d7552;
    ram_cell[     157] = 32'h0;  // 32'hd0003a5d;
    ram_cell[     158] = 32'h0;  // 32'h5806afae;
    ram_cell[     159] = 32'h0;  // 32'hed78ccbc;
    ram_cell[     160] = 32'h0;  // 32'ha07baf85;
    ram_cell[     161] = 32'h0;  // 32'hd13045cd;
    ram_cell[     162] = 32'h0;  // 32'h577680e9;
    ram_cell[     163] = 32'h0;  // 32'hb2165a6d;
    ram_cell[     164] = 32'h0;  // 32'h9e6cc06a;
    ram_cell[     165] = 32'h0;  // 32'hae92affd;
    ram_cell[     166] = 32'h0;  // 32'h133d5ee4;
    ram_cell[     167] = 32'h0;  // 32'h5cb98419;
    ram_cell[     168] = 32'h0;  // 32'h2ef923ee;
    ram_cell[     169] = 32'h0;  // 32'h2843caa9;
    ram_cell[     170] = 32'h0;  // 32'h8eda4caf;
    ram_cell[     171] = 32'h0;  // 32'hf3581bc3;
    ram_cell[     172] = 32'h0;  // 32'h805a7161;
    ram_cell[     173] = 32'h0;  // 32'h63946085;
    ram_cell[     174] = 32'h0;  // 32'hd05e3e68;
    ram_cell[     175] = 32'h0;  // 32'hb65d7b6b;
    ram_cell[     176] = 32'h0;  // 32'h4427120d;
    ram_cell[     177] = 32'h0;  // 32'h20004987;
    ram_cell[     178] = 32'h0;  // 32'he7919a6e;
    ram_cell[     179] = 32'h0;  // 32'h225e5fb7;
    ram_cell[     180] = 32'h0;  // 32'h5e98fc67;
    ram_cell[     181] = 32'h0;  // 32'h3aa27e15;
    ram_cell[     182] = 32'h0;  // 32'hc0184ab3;
    ram_cell[     183] = 32'h0;  // 32'h00f97c24;
    ram_cell[     184] = 32'h0;  // 32'h1538aeae;
    ram_cell[     185] = 32'h0;  // 32'h2dedcdcf;
    ram_cell[     186] = 32'h0;  // 32'h4fedbcda;
    ram_cell[     187] = 32'h0;  // 32'hb0b5137e;
    ram_cell[     188] = 32'h0;  // 32'h9ab55edf;
    ram_cell[     189] = 32'h0;  // 32'h7fad22fa;
    ram_cell[     190] = 32'h0;  // 32'h3790d06f;
    ram_cell[     191] = 32'h0;  // 32'hac33aae2;
    ram_cell[     192] = 32'h0;  // 32'h0ca113fa;
    ram_cell[     193] = 32'h0;  // 32'had07ed64;
    ram_cell[     194] = 32'h0;  // 32'h0f0ab9d1;
    ram_cell[     195] = 32'h0;  // 32'hf0903331;
    ram_cell[     196] = 32'h0;  // 32'hc5e2ea0d;
    ram_cell[     197] = 32'h0;  // 32'hcc978735;
    ram_cell[     198] = 32'h0;  // 32'h666c0d57;
    ram_cell[     199] = 32'h0;  // 32'h00e5c61e;
    ram_cell[     200] = 32'h0;  // 32'h0299cb8e;
    ram_cell[     201] = 32'h0;  // 32'h7216f83c;
    ram_cell[     202] = 32'h0;  // 32'hc4cce8ac;
    ram_cell[     203] = 32'h0;  // 32'h19792e2c;
    ram_cell[     204] = 32'h0;  // 32'he43bc765;
    ram_cell[     205] = 32'h0;  // 32'h1e47be19;
    ram_cell[     206] = 32'h0;  // 32'h9af804bc;
    ram_cell[     207] = 32'h0;  // 32'h9064de35;
    ram_cell[     208] = 32'h0;  // 32'hfe732452;
    ram_cell[     209] = 32'h0;  // 32'h9912e418;
    ram_cell[     210] = 32'h0;  // 32'h4d780995;
    ram_cell[     211] = 32'h0;  // 32'h5e862a9a;
    ram_cell[     212] = 32'h0;  // 32'h06dc0b8f;
    ram_cell[     213] = 32'h0;  // 32'hb9fc180f;
    ram_cell[     214] = 32'h0;  // 32'h6685a7e9;
    ram_cell[     215] = 32'h0;  // 32'h0d9435a8;
    ram_cell[     216] = 32'h0;  // 32'h89d44b62;
    ram_cell[     217] = 32'h0;  // 32'h89a3abd2;
    ram_cell[     218] = 32'h0;  // 32'ha9f4ee48;
    ram_cell[     219] = 32'h0;  // 32'hd113b5b2;
    ram_cell[     220] = 32'h0;  // 32'he141133b;
    ram_cell[     221] = 32'h0;  // 32'hed7189ec;
    ram_cell[     222] = 32'h0;  // 32'h6b36ba60;
    ram_cell[     223] = 32'h0;  // 32'h47210850;
    ram_cell[     224] = 32'h0;  // 32'h323fc389;
    ram_cell[     225] = 32'h0;  // 32'h88ce4aa9;
    ram_cell[     226] = 32'h0;  // 32'hc5c07826;
    ram_cell[     227] = 32'h0;  // 32'hebd064bb;
    ram_cell[     228] = 32'h0;  // 32'h01356236;
    ram_cell[     229] = 32'h0;  // 32'ha562de04;
    ram_cell[     230] = 32'h0;  // 32'h2eb25119;
    ram_cell[     231] = 32'h0;  // 32'h7678d925;
    ram_cell[     232] = 32'h0;  // 32'h9dc8d842;
    ram_cell[     233] = 32'h0;  // 32'hfd3c9b03;
    ram_cell[     234] = 32'h0;  // 32'ha5a53feb;
    ram_cell[     235] = 32'h0;  // 32'ha8c3d8eb;
    ram_cell[     236] = 32'h0;  // 32'h2632e32f;
    ram_cell[     237] = 32'h0;  // 32'he1630232;
    ram_cell[     238] = 32'h0;  // 32'h1dad78fb;
    ram_cell[     239] = 32'h0;  // 32'ha3d20132;
    ram_cell[     240] = 32'h0;  // 32'h721c24a2;
    ram_cell[     241] = 32'h0;  // 32'h960b400e;
    ram_cell[     242] = 32'h0;  // 32'h882f635f;
    ram_cell[     243] = 32'h0;  // 32'h3fb3c0c1;
    ram_cell[     244] = 32'h0;  // 32'h2d7e24c0;
    ram_cell[     245] = 32'h0;  // 32'hc1cef052;
    ram_cell[     246] = 32'h0;  // 32'hfd14f573;
    ram_cell[     247] = 32'h0;  // 32'hd84b674f;
    ram_cell[     248] = 32'h0;  // 32'h62b96728;
    ram_cell[     249] = 32'h0;  // 32'hec99c056;
    ram_cell[     250] = 32'h0;  // 32'h4b528d8c;
    ram_cell[     251] = 32'h0;  // 32'hb1546834;
    ram_cell[     252] = 32'h0;  // 32'h3a2d261a;
    ram_cell[     253] = 32'h0;  // 32'h74afa007;
    ram_cell[     254] = 32'h0;  // 32'h385977e7;
    ram_cell[     255] = 32'h0;  // 32'h026de258;
    // src matrix A
    ram_cell[     256] = 32'h67d8698f;
    ram_cell[     257] = 32'h8c610bcd;
    ram_cell[     258] = 32'h19c31271;
    ram_cell[     259] = 32'h01319e70;
    ram_cell[     260] = 32'h75726570;
    ram_cell[     261] = 32'hcf7242eb;
    ram_cell[     262] = 32'hd8c8dc7e;
    ram_cell[     263] = 32'h061fb4fd;
    ram_cell[     264] = 32'h638dff2d;
    ram_cell[     265] = 32'h91fa4378;
    ram_cell[     266] = 32'h3ecba3a5;
    ram_cell[     267] = 32'hd831b490;
    ram_cell[     268] = 32'ha71bf20f;
    ram_cell[     269] = 32'h69db3bcc;
    ram_cell[     270] = 32'h0c15f397;
    ram_cell[     271] = 32'h9f8c83c4;
    ram_cell[     272] = 32'hacc3c1f2;
    ram_cell[     273] = 32'h2fc9076d;
    ram_cell[     274] = 32'h56aa590e;
    ram_cell[     275] = 32'h0ed45912;
    ram_cell[     276] = 32'h9ee5a817;
    ram_cell[     277] = 32'he7f5ab3b;
    ram_cell[     278] = 32'hf8cc599c;
    ram_cell[     279] = 32'h16d6f4d7;
    ram_cell[     280] = 32'he0ec4b29;
    ram_cell[     281] = 32'h6e4451a4;
    ram_cell[     282] = 32'h716d45a6;
    ram_cell[     283] = 32'h57c8ec28;
    ram_cell[     284] = 32'hf883e01c;
    ram_cell[     285] = 32'hf059b62c;
    ram_cell[     286] = 32'hc5a42bdf;
    ram_cell[     287] = 32'he452668e;
    ram_cell[     288] = 32'hf5f6d84c;
    ram_cell[     289] = 32'h6854d378;
    ram_cell[     290] = 32'he64c55dd;
    ram_cell[     291] = 32'h76ca6254;
    ram_cell[     292] = 32'h70eebbe9;
    ram_cell[     293] = 32'hc8a01dea;
    ram_cell[     294] = 32'he0ed2d64;
    ram_cell[     295] = 32'h7b18bb4a;
    ram_cell[     296] = 32'h2a011dc1;
    ram_cell[     297] = 32'h4ae139e9;
    ram_cell[     298] = 32'h58686830;
    ram_cell[     299] = 32'h5fe3d6d0;
    ram_cell[     300] = 32'h4e77239c;
    ram_cell[     301] = 32'h494f7e33;
    ram_cell[     302] = 32'hf01be2d6;
    ram_cell[     303] = 32'hcc775147;
    ram_cell[     304] = 32'ha1ba8233;
    ram_cell[     305] = 32'h6e097f80;
    ram_cell[     306] = 32'h1f4a81be;
    ram_cell[     307] = 32'h62df4af8;
    ram_cell[     308] = 32'h92370d52;
    ram_cell[     309] = 32'hd213a904;
    ram_cell[     310] = 32'h47ed0b92;
    ram_cell[     311] = 32'h88b1ef57;
    ram_cell[     312] = 32'h50f6c490;
    ram_cell[     313] = 32'h161fba2f;
    ram_cell[     314] = 32'hc4ac7e33;
    ram_cell[     315] = 32'hc1a11315;
    ram_cell[     316] = 32'h0aeaf494;
    ram_cell[     317] = 32'hc7748b0d;
    ram_cell[     318] = 32'hc729c5cf;
    ram_cell[     319] = 32'h271ce229;
    ram_cell[     320] = 32'heee9724d;
    ram_cell[     321] = 32'ha309e1ca;
    ram_cell[     322] = 32'hce2d1c8c;
    ram_cell[     323] = 32'h5a65d46b;
    ram_cell[     324] = 32'h3fb15061;
    ram_cell[     325] = 32'hb214bff3;
    ram_cell[     326] = 32'hc093efbb;
    ram_cell[     327] = 32'hb065aacd;
    ram_cell[     328] = 32'h35bc1942;
    ram_cell[     329] = 32'hb3476408;
    ram_cell[     330] = 32'h63fb4c9b;
    ram_cell[     331] = 32'h92b4825e;
    ram_cell[     332] = 32'h8bc52ab7;
    ram_cell[     333] = 32'h54e794bd;
    ram_cell[     334] = 32'h5e2ac6c7;
    ram_cell[     335] = 32'h10cd7711;
    ram_cell[     336] = 32'h572c1d36;
    ram_cell[     337] = 32'hb3921e4d;
    ram_cell[     338] = 32'h23ff7d7d;
    ram_cell[     339] = 32'hf27f6326;
    ram_cell[     340] = 32'ha3bf777e;
    ram_cell[     341] = 32'h78f96c64;
    ram_cell[     342] = 32'h51c8faa2;
    ram_cell[     343] = 32'hf0067422;
    ram_cell[     344] = 32'h42942dd8;
    ram_cell[     345] = 32'h41126140;
    ram_cell[     346] = 32'ha88dbbc8;
    ram_cell[     347] = 32'hcc5631c9;
    ram_cell[     348] = 32'h14404329;
    ram_cell[     349] = 32'hc965fb86;
    ram_cell[     350] = 32'hb0a0647a;
    ram_cell[     351] = 32'hff364362;
    ram_cell[     352] = 32'h5b840b91;
    ram_cell[     353] = 32'h2e4013f9;
    ram_cell[     354] = 32'hdbca2c70;
    ram_cell[     355] = 32'h8cebbbd0;
    ram_cell[     356] = 32'hc9434d0c;
    ram_cell[     357] = 32'h367eca05;
    ram_cell[     358] = 32'hc4122dcf;
    ram_cell[     359] = 32'h678532a4;
    ram_cell[     360] = 32'ha7e90b1d;
    ram_cell[     361] = 32'h96ed26ff;
    ram_cell[     362] = 32'haf030c63;
    ram_cell[     363] = 32'hd15f3079;
    ram_cell[     364] = 32'hab9121e9;
    ram_cell[     365] = 32'h88a1a762;
    ram_cell[     366] = 32'h761088e4;
    ram_cell[     367] = 32'h592a3a48;
    ram_cell[     368] = 32'h1ed41ea3;
    ram_cell[     369] = 32'h9cd727f8;
    ram_cell[     370] = 32'he35ebc52;
    ram_cell[     371] = 32'h98115589;
    ram_cell[     372] = 32'h7be53967;
    ram_cell[     373] = 32'hec099c90;
    ram_cell[     374] = 32'h86d629b5;
    ram_cell[     375] = 32'h42becd58;
    ram_cell[     376] = 32'h1007ab6c;
    ram_cell[     377] = 32'h37a512cb;
    ram_cell[     378] = 32'h65f817c8;
    ram_cell[     379] = 32'h471d6ba6;
    ram_cell[     380] = 32'he5e03cf5;
    ram_cell[     381] = 32'hb499633c;
    ram_cell[     382] = 32'h7f9240bb;
    ram_cell[     383] = 32'h5c882cde;
    ram_cell[     384] = 32'h488e3f72;
    ram_cell[     385] = 32'h4c0fcbb9;
    ram_cell[     386] = 32'hac1005ce;
    ram_cell[     387] = 32'h2faaf454;
    ram_cell[     388] = 32'hc65d9649;
    ram_cell[     389] = 32'heefc4c5f;
    ram_cell[     390] = 32'h43949eef;
    ram_cell[     391] = 32'h6becd86a;
    ram_cell[     392] = 32'hdd098073;
    ram_cell[     393] = 32'h8f6639bb;
    ram_cell[     394] = 32'hf0de0b7d;
    ram_cell[     395] = 32'h505b26e4;
    ram_cell[     396] = 32'he5b151d0;
    ram_cell[     397] = 32'h5d08f36e;
    ram_cell[     398] = 32'h348ab947;
    ram_cell[     399] = 32'h206865bf;
    ram_cell[     400] = 32'h88357a1e;
    ram_cell[     401] = 32'h7575f860;
    ram_cell[     402] = 32'h04c0902b;
    ram_cell[     403] = 32'h569809e4;
    ram_cell[     404] = 32'h27faf234;
    ram_cell[     405] = 32'h0d275d4e;
    ram_cell[     406] = 32'h77592712;
    ram_cell[     407] = 32'hf67df140;
    ram_cell[     408] = 32'hf1a468cc;
    ram_cell[     409] = 32'h447c87c6;
    ram_cell[     410] = 32'ha64c2902;
    ram_cell[     411] = 32'h7b26b6c5;
    ram_cell[     412] = 32'hf765005f;
    ram_cell[     413] = 32'h74596958;
    ram_cell[     414] = 32'ha93327e8;
    ram_cell[     415] = 32'h7726301a;
    ram_cell[     416] = 32'hccf47dff;
    ram_cell[     417] = 32'h791ab941;
    ram_cell[     418] = 32'h482dddf4;
    ram_cell[     419] = 32'hdeea602b;
    ram_cell[     420] = 32'h9ecb7331;
    ram_cell[     421] = 32'h0a83b4a2;
    ram_cell[     422] = 32'h309d6a9e;
    ram_cell[     423] = 32'h07210c69;
    ram_cell[     424] = 32'h94b51512;
    ram_cell[     425] = 32'h5ce6933b;
    ram_cell[     426] = 32'h5495363e;
    ram_cell[     427] = 32'he01a32d2;
    ram_cell[     428] = 32'h95f01489;
    ram_cell[     429] = 32'ha779f64f;
    ram_cell[     430] = 32'h8e3c3655;
    ram_cell[     431] = 32'h40a482c3;
    ram_cell[     432] = 32'h359c7995;
    ram_cell[     433] = 32'h2dac5e11;
    ram_cell[     434] = 32'h1fc8bbb3;
    ram_cell[     435] = 32'h5b40cca4;
    ram_cell[     436] = 32'hd6100397;
    ram_cell[     437] = 32'h1a8e41e9;
    ram_cell[     438] = 32'h16a738bc;
    ram_cell[     439] = 32'h45194550;
    ram_cell[     440] = 32'hef23dd21;
    ram_cell[     441] = 32'hc985c999;
    ram_cell[     442] = 32'h475798b6;
    ram_cell[     443] = 32'h99061f65;
    ram_cell[     444] = 32'h6e56f2a2;
    ram_cell[     445] = 32'h84caeb77;
    ram_cell[     446] = 32'hce2850e0;
    ram_cell[     447] = 32'h22496a98;
    ram_cell[     448] = 32'hcacbe4e4;
    ram_cell[     449] = 32'hb7a7ac61;
    ram_cell[     450] = 32'h19a9312e;
    ram_cell[     451] = 32'h295324d3;
    ram_cell[     452] = 32'h00515513;
    ram_cell[     453] = 32'h1b2bdea6;
    ram_cell[     454] = 32'h986f2ecf;
    ram_cell[     455] = 32'h134bbe72;
    ram_cell[     456] = 32'h2478ee3c;
    ram_cell[     457] = 32'h52b84505;
    ram_cell[     458] = 32'h1d15dfc2;
    ram_cell[     459] = 32'he9d78654;
    ram_cell[     460] = 32'h26760ba3;
    ram_cell[     461] = 32'h3fd5c422;
    ram_cell[     462] = 32'h6ef65798;
    ram_cell[     463] = 32'haaf69cce;
    ram_cell[     464] = 32'h7738536c;
    ram_cell[     465] = 32'ha2a82a7a;
    ram_cell[     466] = 32'h7a3a2aa9;
    ram_cell[     467] = 32'h0b4ec007;
    ram_cell[     468] = 32'hb5573a1d;
    ram_cell[     469] = 32'hd0dc8ab7;
    ram_cell[     470] = 32'h4b733a9a;
    ram_cell[     471] = 32'h933313c4;
    ram_cell[     472] = 32'h62205d38;
    ram_cell[     473] = 32'h4726e417;
    ram_cell[     474] = 32'hb86e3365;
    ram_cell[     475] = 32'h85e7513d;
    ram_cell[     476] = 32'h2903fe7f;
    ram_cell[     477] = 32'h0ee40d72;
    ram_cell[     478] = 32'h7697ad9c;
    ram_cell[     479] = 32'h24efcd6a;
    ram_cell[     480] = 32'ha3a32460;
    ram_cell[     481] = 32'h876de780;
    ram_cell[     482] = 32'hf3383aa2;
    ram_cell[     483] = 32'h8fdd9ce3;
    ram_cell[     484] = 32'h877b7f9e;
    ram_cell[     485] = 32'hc6608297;
    ram_cell[     486] = 32'hfcd0aefc;
    ram_cell[     487] = 32'he2bdb75b;
    ram_cell[     488] = 32'h701da6a1;
    ram_cell[     489] = 32'h262bd0a0;
    ram_cell[     490] = 32'h21aca32c;
    ram_cell[     491] = 32'h70a3a005;
    ram_cell[     492] = 32'he202d04a;
    ram_cell[     493] = 32'h3a220663;
    ram_cell[     494] = 32'ha2758f14;
    ram_cell[     495] = 32'h71548279;
    ram_cell[     496] = 32'hec408e79;
    ram_cell[     497] = 32'he4b5879b;
    ram_cell[     498] = 32'h0807488c;
    ram_cell[     499] = 32'h14dbefb9;
    ram_cell[     500] = 32'h5dd6b844;
    ram_cell[     501] = 32'h8da7497a;
    ram_cell[     502] = 32'hf9b38157;
    ram_cell[     503] = 32'hde377702;
    ram_cell[     504] = 32'hd4acd99b;
    ram_cell[     505] = 32'h14cee8cf;
    ram_cell[     506] = 32'hac447fc5;
    ram_cell[     507] = 32'h3bb6a131;
    ram_cell[     508] = 32'hf89d1e30;
    ram_cell[     509] = 32'h35a92b57;
    ram_cell[     510] = 32'ha9316031;
    ram_cell[     511] = 32'h5bfc4f07;
    // src matrix B
    ram_cell[     512] = 32'h1f45a398;
    ram_cell[     513] = 32'h57bf5d68;
    ram_cell[     514] = 32'h6e830ed6;
    ram_cell[     515] = 32'h42858764;
    ram_cell[     516] = 32'h42dc241a;
    ram_cell[     517] = 32'hd9b5abd1;
    ram_cell[     518] = 32'h33544f33;
    ram_cell[     519] = 32'h69c9ae7c;
    ram_cell[     520] = 32'h03343fef;
    ram_cell[     521] = 32'h564b7a8f;
    ram_cell[     522] = 32'h21f69f72;
    ram_cell[     523] = 32'h164421e7;
    ram_cell[     524] = 32'h41d65f02;
    ram_cell[     525] = 32'hb7201540;
    ram_cell[     526] = 32'h03d476b1;
    ram_cell[     527] = 32'hd8513938;
    ram_cell[     528] = 32'had693a1e;
    ram_cell[     529] = 32'h57423a0e;
    ram_cell[     530] = 32'hdf5c8ed4;
    ram_cell[     531] = 32'h44e6067f;
    ram_cell[     532] = 32'h0de1908d;
    ram_cell[     533] = 32'h0daf9884;
    ram_cell[     534] = 32'hd540f4c9;
    ram_cell[     535] = 32'h96290e6a;
    ram_cell[     536] = 32'h2a2ac124;
    ram_cell[     537] = 32'hb44b6099;
    ram_cell[     538] = 32'hf3b54388;
    ram_cell[     539] = 32'h26415dd7;
    ram_cell[     540] = 32'hab94abb1;
    ram_cell[     541] = 32'h04f0c498;
    ram_cell[     542] = 32'hcc988373;
    ram_cell[     543] = 32'h3405a855;
    ram_cell[     544] = 32'h9783c322;
    ram_cell[     545] = 32'hee028d1e;
    ram_cell[     546] = 32'h57cba0f1;
    ram_cell[     547] = 32'hbba73170;
    ram_cell[     548] = 32'h2dad5b05;
    ram_cell[     549] = 32'hfd2b9983;
    ram_cell[     550] = 32'hb736d670;
    ram_cell[     551] = 32'hbe29bfbf;
    ram_cell[     552] = 32'h38eaafde;
    ram_cell[     553] = 32'hea4a8466;
    ram_cell[     554] = 32'h8adae90e;
    ram_cell[     555] = 32'h81f85c27;
    ram_cell[     556] = 32'h686beb03;
    ram_cell[     557] = 32'h88c015d1;
    ram_cell[     558] = 32'h3c162f2c;
    ram_cell[     559] = 32'h167d0174;
    ram_cell[     560] = 32'h2ccc3211;
    ram_cell[     561] = 32'hcbd3ebd9;
    ram_cell[     562] = 32'hc04c058e;
    ram_cell[     563] = 32'h43c9acb1;
    ram_cell[     564] = 32'h01f3b5b2;
    ram_cell[     565] = 32'hcc22277f;
    ram_cell[     566] = 32'h8fbac4eb;
    ram_cell[     567] = 32'hffa34e39;
    ram_cell[     568] = 32'h3ee2bb13;
    ram_cell[     569] = 32'hbdffc1bb;
    ram_cell[     570] = 32'hc8d8e37f;
    ram_cell[     571] = 32'h5bd4094a;
    ram_cell[     572] = 32'h77d31335;
    ram_cell[     573] = 32'h9093dd55;
    ram_cell[     574] = 32'h36daeebf;
    ram_cell[     575] = 32'h7ef51610;
    ram_cell[     576] = 32'ha0b5cd94;
    ram_cell[     577] = 32'h83e5a158;
    ram_cell[     578] = 32'h613c5e6b;
    ram_cell[     579] = 32'h6fe61445;
    ram_cell[     580] = 32'hcd30d4cd;
    ram_cell[     581] = 32'h47176ca1;
    ram_cell[     582] = 32'ha17d701f;
    ram_cell[     583] = 32'h04d0e4cd;
    ram_cell[     584] = 32'hb963addf;
    ram_cell[     585] = 32'hd862ec76;
    ram_cell[     586] = 32'h201bd7b2;
    ram_cell[     587] = 32'h6d9b99c1;
    ram_cell[     588] = 32'hf828c73e;
    ram_cell[     589] = 32'ha102c080;
    ram_cell[     590] = 32'h88902d0e;
    ram_cell[     591] = 32'h1752e9b4;
    ram_cell[     592] = 32'hd89baf0a;
    ram_cell[     593] = 32'h4d94aa75;
    ram_cell[     594] = 32'hd116dddf;
    ram_cell[     595] = 32'hf7a07ae7;
    ram_cell[     596] = 32'h71326ca0;
    ram_cell[     597] = 32'h9ed0fe3e;
    ram_cell[     598] = 32'hac115ae8;
    ram_cell[     599] = 32'h4d7b4a28;
    ram_cell[     600] = 32'h04671e9b;
    ram_cell[     601] = 32'ha4fce8bc;
    ram_cell[     602] = 32'hb88989ff;
    ram_cell[     603] = 32'hf67b2945;
    ram_cell[     604] = 32'h04babb6e;
    ram_cell[     605] = 32'heb5f39a5;
    ram_cell[     606] = 32'hac603dd3;
    ram_cell[     607] = 32'h22afed6f;
    ram_cell[     608] = 32'h205393fe;
    ram_cell[     609] = 32'h4894e651;
    ram_cell[     610] = 32'h377f2619;
    ram_cell[     611] = 32'h34d01769;
    ram_cell[     612] = 32'h1b095dff;
    ram_cell[     613] = 32'hd47b7f5d;
    ram_cell[     614] = 32'haa2b8d9a;
    ram_cell[     615] = 32'h0d9ff01d;
    ram_cell[     616] = 32'h319917af;
    ram_cell[     617] = 32'h787d35d6;
    ram_cell[     618] = 32'h456c5ffc;
    ram_cell[     619] = 32'hc9ab36fc;
    ram_cell[     620] = 32'hdb847dae;
    ram_cell[     621] = 32'hdf925627;
    ram_cell[     622] = 32'h1431213c;
    ram_cell[     623] = 32'h8489e552;
    ram_cell[     624] = 32'h90905fd2;
    ram_cell[     625] = 32'hb9b5b86a;
    ram_cell[     626] = 32'ha23926c6;
    ram_cell[     627] = 32'hac82bcbf;
    ram_cell[     628] = 32'hb4cfa197;
    ram_cell[     629] = 32'h11c38482;
    ram_cell[     630] = 32'h31e9a51e;
    ram_cell[     631] = 32'hd500c7fb;
    ram_cell[     632] = 32'hc71586d0;
    ram_cell[     633] = 32'hefd3d750;
    ram_cell[     634] = 32'hf00faea0;
    ram_cell[     635] = 32'h866bc2f6;
    ram_cell[     636] = 32'h2fb70004;
    ram_cell[     637] = 32'hfb60c440;
    ram_cell[     638] = 32'he30d9ddc;
    ram_cell[     639] = 32'h54ceb06a;
    ram_cell[     640] = 32'h0bbc320a;
    ram_cell[     641] = 32'h16fc0b87;
    ram_cell[     642] = 32'h3ddf0c16;
    ram_cell[     643] = 32'h3fd1e8b2;
    ram_cell[     644] = 32'h32898950;
    ram_cell[     645] = 32'h4b02d7df;
    ram_cell[     646] = 32'hf2de3066;
    ram_cell[     647] = 32'hbc73c353;
    ram_cell[     648] = 32'h13211bf9;
    ram_cell[     649] = 32'h80ea5afc;
    ram_cell[     650] = 32'h2a991ce1;
    ram_cell[     651] = 32'hc036e49e;
    ram_cell[     652] = 32'h9f33a052;
    ram_cell[     653] = 32'hf6059075;
    ram_cell[     654] = 32'h605a8c51;
    ram_cell[     655] = 32'h7f205a1a;
    ram_cell[     656] = 32'h0cb461e6;
    ram_cell[     657] = 32'h8c6a84e3;
    ram_cell[     658] = 32'hfdb361fa;
    ram_cell[     659] = 32'he141ef60;
    ram_cell[     660] = 32'habc58f74;
    ram_cell[     661] = 32'hb0a3d37c;
    ram_cell[     662] = 32'h014b4a6f;
    ram_cell[     663] = 32'h85d8ba7d;
    ram_cell[     664] = 32'h508956f6;
    ram_cell[     665] = 32'h847afaf8;
    ram_cell[     666] = 32'hea021e42;
    ram_cell[     667] = 32'he904d5ad;
    ram_cell[     668] = 32'ha4184d68;
    ram_cell[     669] = 32'h0a1aa713;
    ram_cell[     670] = 32'h98005098;
    ram_cell[     671] = 32'h051e57d4;
    ram_cell[     672] = 32'h88b6408b;
    ram_cell[     673] = 32'h55d3b824;
    ram_cell[     674] = 32'hbcb77e74;
    ram_cell[     675] = 32'h0e32935d;
    ram_cell[     676] = 32'h63c4ed08;
    ram_cell[     677] = 32'h79cfd126;
    ram_cell[     678] = 32'h6f78d0a0;
    ram_cell[     679] = 32'h4ce2e6e8;
    ram_cell[     680] = 32'h195e02d5;
    ram_cell[     681] = 32'hff2c054b;
    ram_cell[     682] = 32'heab69c65;
    ram_cell[     683] = 32'h121bd723;
    ram_cell[     684] = 32'h3eb2bf0a;
    ram_cell[     685] = 32'h20045318;
    ram_cell[     686] = 32'h85a98680;
    ram_cell[     687] = 32'h23b1e949;
    ram_cell[     688] = 32'h6bcfc8b3;
    ram_cell[     689] = 32'he44aa120;
    ram_cell[     690] = 32'h70ee7ff5;
    ram_cell[     691] = 32'hda8ef655;
    ram_cell[     692] = 32'hd264e3dd;
    ram_cell[     693] = 32'h1701f7d2;
    ram_cell[     694] = 32'ha18c04fb;
    ram_cell[     695] = 32'hacc3dbb2;
    ram_cell[     696] = 32'h185999bd;
    ram_cell[     697] = 32'h0bc8c16a;
    ram_cell[     698] = 32'h202af294;
    ram_cell[     699] = 32'h27a95688;
    ram_cell[     700] = 32'h50131712;
    ram_cell[     701] = 32'hc98bffec;
    ram_cell[     702] = 32'h2aba8362;
    ram_cell[     703] = 32'ha46120ca;
    ram_cell[     704] = 32'hec68970d;
    ram_cell[     705] = 32'h68a2d137;
    ram_cell[     706] = 32'h323c0ab3;
    ram_cell[     707] = 32'h5d64c667;
    ram_cell[     708] = 32'h0f9ce166;
    ram_cell[     709] = 32'he05ca8c6;
    ram_cell[     710] = 32'h05c5e96f;
    ram_cell[     711] = 32'h6d2ab47a;
    ram_cell[     712] = 32'h99479a5f;
    ram_cell[     713] = 32'h3c2994aa;
    ram_cell[     714] = 32'hb28d2b97;
    ram_cell[     715] = 32'h15ed2c5f;
    ram_cell[     716] = 32'h54b0af91;
    ram_cell[     717] = 32'h8b183096;
    ram_cell[     718] = 32'ha1b7f59c;
    ram_cell[     719] = 32'hee907e92;
    ram_cell[     720] = 32'h4246b360;
    ram_cell[     721] = 32'h5d611844;
    ram_cell[     722] = 32'h18e0ef46;
    ram_cell[     723] = 32'h7eeaeb61;
    ram_cell[     724] = 32'h476fefad;
    ram_cell[     725] = 32'h4b579daf;
    ram_cell[     726] = 32'hd6c1e4d6;
    ram_cell[     727] = 32'h517ab428;
    ram_cell[     728] = 32'h051f8a47;
    ram_cell[     729] = 32'h1545ecc1;
    ram_cell[     730] = 32'h5f8ce6d2;
    ram_cell[     731] = 32'h5a72b7aa;
    ram_cell[     732] = 32'h13934cc3;
    ram_cell[     733] = 32'h1753d480;
    ram_cell[     734] = 32'h148a9e0d;
    ram_cell[     735] = 32'hdcc41aa2;
    ram_cell[     736] = 32'hf1da2eb2;
    ram_cell[     737] = 32'h414ae618;
    ram_cell[     738] = 32'hd8b80ec7;
    ram_cell[     739] = 32'h4c9da62b;
    ram_cell[     740] = 32'hd4d524a1;
    ram_cell[     741] = 32'hd3c1f1f0;
    ram_cell[     742] = 32'h8974369b;
    ram_cell[     743] = 32'h863b1f8d;
    ram_cell[     744] = 32'h680bf9d8;
    ram_cell[     745] = 32'h3df3e6cc;
    ram_cell[     746] = 32'h125305cd;
    ram_cell[     747] = 32'h0ef23fa8;
    ram_cell[     748] = 32'hd262f4a0;
    ram_cell[     749] = 32'hd4f40ab8;
    ram_cell[     750] = 32'h238f19a1;
    ram_cell[     751] = 32'hd12b67c3;
    ram_cell[     752] = 32'h41e3eae7;
    ram_cell[     753] = 32'hf94ea92e;
    ram_cell[     754] = 32'h97ae03ba;
    ram_cell[     755] = 32'hf243749a;
    ram_cell[     756] = 32'h12fe7deb;
    ram_cell[     757] = 32'hcd717b35;
    ram_cell[     758] = 32'h35cade2f;
    ram_cell[     759] = 32'hbcd247cc;
    ram_cell[     760] = 32'haebb8a49;
    ram_cell[     761] = 32'hb59ed75b;
    ram_cell[     762] = 32'h1cf086f6;
    ram_cell[     763] = 32'hee2286ac;
    ram_cell[     764] = 32'hc1bfe057;
    ram_cell[     765] = 32'hded0780b;
    ram_cell[     766] = 32'h1ae9f25d;
    ram_cell[     767] = 32'h8453a717;
    
end

endmodule

